-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"880b0b0b",
     1 => x"0b81e004",
     2 => x"8804ff0d",
     3 => x"80040000",
     4 => x"80e0040b",
     5 => x"80f5040b",
     6 => x"81a2040b",
     7 => x"81b70404",
     8 => x"0b0b0bbc",
     9 => x"8c080b0b",
    10 => x"0bbc9008",
    11 => x"0b0b0bbc",
    12 => x"94080b0b",
    13 => x"0b80cc08",
    14 => x"2d0b0b0b",
    15 => x"bc940c0b",
    16 => x"0b0bbc90",
    17 => x"0c0b0b0b",
    18 => x"bc8c0c04",
    19 => x"0000001f",
    20 => x"00ffffff",
    21 => x"ff00ffff",
    22 => x"ffff00ff",
    23 => x"ffffff00",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fd06",
    30 => x"0883ffff",
    31 => x"73830609",
    32 => x"81058205",
    33 => x"832b2b09",
    34 => x"067383ff",
    35 => x"ff067383",
    36 => x"06098105",
    37 => x"8205832b",
    38 => x"0b2b0772",
    39 => x"fc060c51",
    40 => x"510471fc",
    41 => x"06087283",
    42 => x"06098105",
    43 => x"83051010",
    44 => x"102a81ff",
    45 => x"06520471",
    46 => x"fc06080b",
    47 => x"0b0b80d0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bc8c7080",
    57 => x"c6cc278e",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"0b0b0b81",
    61 => x"e2048851",
    62 => x"8fc30402",
    63 => x"fc050df8",
    64 => x"80518f0b",
    65 => x"bc9c0c9f",
    66 => x"0bbca00c",
    67 => x"a0717081",
    68 => x"055334bc",
    69 => x"a008ff05",
    70 => x"bca00cbc",
    71 => x"a0088025",
    72 => x"eb38bc9c",
    73 => x"08ff05bc",
    74 => x"9c0cbc9c",
    75 => x"088025d7",
    76 => x"38028405",
    77 => x"0d0402f0",
    78 => x"050df880",
    79 => x"53f8a054",
    80 => x"83bf5273",
    81 => x"70810555",
    82 => x"33517073",
    83 => x"70810555",
    84 => x"34ff1252",
    85 => x"718025eb",
    86 => x"38fbc053",
    87 => x"9f52a073",
    88 => x"70810555",
    89 => x"34ff1252",
    90 => x"718025f2",
    91 => x"38029005",
    92 => x"0d0402f4",
    93 => x"050d7453",
    94 => x"8e0bbc9c",
    95 => x"08258f38",
    96 => x"82b62dbc",
    97 => x"9c08ff05",
    98 => x"bc9c0c82",
    99 => x"f804bc9c",
   100 => x"08bca008",
   101 => x"5351728a",
   102 => x"2e098106",
   103 => x"b7387151",
   104 => x"719f24a0",
   105 => x"38bc9c08",
   106 => x"a02911f8",
   107 => x"80115151",
   108 => x"a07134bc",
   109 => x"a0088105",
   110 => x"bca00cbc",
   111 => x"a008519f",
   112 => x"7125e238",
   113 => x"800bbca0",
   114 => x"0cbc9c08",
   115 => x"8105bc9c",
   116 => x"0c83e804",
   117 => x"70a02912",
   118 => x"f8801151",
   119 => x"51727134",
   120 => x"bca00881",
   121 => x"05bca00c",
   122 => x"bca008a0",
   123 => x"2e098106",
   124 => x"8e38800b",
   125 => x"bca00cbc",
   126 => x"9c088105",
   127 => x"bc9c0c02",
   128 => x"8c050d04",
   129 => x"02e8050d",
   130 => x"77795656",
   131 => x"880bfc16",
   132 => x"77712c8f",
   133 => x"06545254",
   134 => x"80537272",
   135 => x"25953871",
   136 => x"53fbe014",
   137 => x"51877134",
   138 => x"8114ff14",
   139 => x"545472f1",
   140 => x"387153f9",
   141 => x"1576712c",
   142 => x"87065351",
   143 => x"71802e8b",
   144 => x"38fbe014",
   145 => x"51717134",
   146 => x"81145472",
   147 => x"8e249538",
   148 => x"8f733153",
   149 => x"fbe01451",
   150 => x"a0713481",
   151 => x"14ff1454",
   152 => x"5472f138",
   153 => x"0298050d",
   154 => x"0402ec05",
   155 => x"0d800bbc",
   156 => x"a40cf68c",
   157 => x"08f69008",
   158 => x"71882c56",
   159 => x"5481ff06",
   160 => x"52737225",
   161 => x"88387154",
   162 => x"820bbca4",
   163 => x"0c72882c",
   164 => x"7381ff06",
   165 => x"54557473",
   166 => x"258b3872",
   167 => x"bca40884",
   168 => x"07bca40c",
   169 => x"5573842b",
   170 => x"87e87125",
   171 => x"83713170",
   172 => x"0b0b0bb8",
   173 => x"f80c8171",
   174 => x"2bf6880c",
   175 => x"fea413ff",
   176 => x"122c7888",
   177 => x"29ff9405",
   178 => x"70812cbc",
   179 => x"a4085258",
   180 => x"52555152",
   181 => x"5476802e",
   182 => x"85387081",
   183 => x"075170f6",
   184 => x"940c7109",
   185 => x"8105f680",
   186 => x"0c720981",
   187 => x"05f6840c",
   188 => x"0294050d",
   189 => x"0402f405",
   190 => x"0d745372",
   191 => x"70810554",
   192 => x"33527180",
   193 => x"2e893871",
   194 => x"5182f22d",
   195 => x"85fb0402",
   196 => x"8c050d04",
   197 => x"02f4050d",
   198 => x"74708206",
   199 => x"80c6b00c",
   200 => x"b9947181",
   201 => x"06545451",
   202 => x"71881434",
   203 => x"70822a70",
   204 => x"81065151",
   205 => x"70a01434",
   206 => x"70bc8c0c",
   207 => x"028c050d",
   208 => x"0402f805",
   209 => x"0d0b0b0b",
   210 => x"b79052bc",
   211 => x"a8519b83",
   212 => x"2dbc8c08",
   213 => x"802e9d38",
   214 => x"bfc452bc",
   215 => x"a8519dba",
   216 => x"2dbfc408",
   217 => x"bcb40cbf",
   218 => x"c408fec0",
   219 => x"0cbfc408",
   220 => x"5186942d",
   221 => x"0288050d",
   222 => x"0402f005",
   223 => x"0d805192",
   224 => x"812d0b0b",
   225 => x"0bb79052",
   226 => x"bca8519b",
   227 => x"832dbc8c",
   228 => x"08802ea5",
   229 => x"38bcb408",
   230 => x"bfc40cbf",
   231 => x"c85480fd",
   232 => x"53807470",
   233 => x"8405560c",
   234 => x"ff135372",
   235 => x"8025f238",
   236 => x"bfc452bc",
   237 => x"a8519de3",
   238 => x"2d029005",
   239 => x"0d0402d4",
   240 => x"050dbcb4",
   241 => x"08fec00c",
   242 => x"810bfec4",
   243 => x"0c840bfe",
   244 => x"c40c7c52",
   245 => x"bca8519b",
   246 => x"832dbc8c",
   247 => x"0853bc8c",
   248 => x"08802e81",
   249 => x"cc38bcac",
   250 => x"0856800b",
   251 => x"ff175859",
   252 => x"76792e8b",
   253 => x"38811977",
   254 => x"812a5859",
   255 => x"76f738f7",
   256 => x"19769fff",
   257 => x"06545972",
   258 => x"802e8b38",
   259 => x"fc8016bc",
   260 => x"a852569d",
   261 => x"8c2d75b0",
   262 => x"80802e09",
   263 => x"81068938",
   264 => x"820bfedc",
   265 => x"0c88bf04",
   266 => x"75988080",
   267 => x"2e098106",
   268 => x"8938810b",
   269 => x"fedc0c88",
   270 => x"bf04800b",
   271 => x"fedc0c81",
   272 => x"5b807625",
   273 => x"80e93878",
   274 => x"52765184",
   275 => x"842dbfc4",
   276 => x"52bca851",
   277 => x"9dba2dbc",
   278 => x"8c08802e",
   279 => x"bb38bfc4",
   280 => x"5a83fc58",
   281 => x"79708405",
   282 => x"5b087083",
   283 => x"fe800671",
   284 => x"882b83fe",
   285 => x"80067188",
   286 => x"2a077288",
   287 => x"2a83fe80",
   288 => x"0673982a",
   289 => x"07fec80c",
   290 => x"fec80c56",
   291 => x"fc195953",
   292 => x"778025d0",
   293 => x"38899f04",
   294 => x"bc8c085b",
   295 => x"848056bc",
   296 => x"a8519d8c",
   297 => x"2dfc8016",
   298 => x"81185856",
   299 => x"88c1047a",
   300 => x"5372bc8c",
   301 => x"0c02ac05",
   302 => x"0d0402fc",
   303 => x"050daadf",
   304 => x"2dfec451",
   305 => x"81710c82",
   306 => x"710c0284",
   307 => x"050d0402",
   308 => x"f4050d74",
   309 => x"76785354",
   310 => x"52807125",
   311 => x"93387270",
   312 => x"81055433",
   313 => x"72708105",
   314 => x"5434ff11",
   315 => x"5170ef38",
   316 => x"80723402",
   317 => x"8c050d04",
   318 => x"02e8050d",
   319 => x"77568070",
   320 => x"56547376",
   321 => x"24b33880",
   322 => x"c5d40874",
   323 => x"2eab3873",
   324 => x"5199892d",
   325 => x"bc8c08bc",
   326 => x"8c080981",
   327 => x"0570bc8c",
   328 => x"08079f2a",
   329 => x"77058117",
   330 => x"57575353",
   331 => x"74762489",
   332 => x"3880c5d4",
   333 => x"087426d7",
   334 => x"3872bc8c",
   335 => x"0c029805",
   336 => x"0d0402f4",
   337 => x"050dbbb8",
   338 => x"08155189",
   339 => x"f82dbc8c",
   340 => x"08802e95",
   341 => x"388b53bc",
   342 => x"8c085280",
   343 => x"c3c45189",
   344 => x"cf2d80c3",
   345 => x"c45187be",
   346 => x"2db8fc51",
   347 => x"acbd2daa",
   348 => x"df2d8051",
   349 => x"84e92d02",
   350 => x"8c050d04",
   351 => x"02dc050d",
   352 => x"80705a55",
   353 => x"74bbb808",
   354 => x"25b13880",
   355 => x"c5d40875",
   356 => x"2ea93878",
   357 => x"5199892d",
   358 => x"bc8c0809",
   359 => x"810570bc",
   360 => x"8c08079f",
   361 => x"2a760581",
   362 => x"1b5b5654",
   363 => x"74bbb808",
   364 => x"25893880",
   365 => x"c5d40879",
   366 => x"26d93880",
   367 => x"557880c5",
   368 => x"d4082781",
   369 => x"c5387851",
   370 => x"99892dbc",
   371 => x"8c08802e",
   372 => x"819c38bc",
   373 => x"8c088b05",
   374 => x"3370842a",
   375 => x"70810677",
   376 => x"1078842b",
   377 => x"80c3c433",
   378 => x"5c5c5351",
   379 => x"55567380",
   380 => x"2e80c338",
   381 => x"7416822b",
   382 => x"8dab0bba",
   383 => x"8c120c54",
   384 => x"77753110",
   385 => x"bcbc1155",
   386 => x"56907470",
   387 => x"81055634",
   388 => x"a0743476",
   389 => x"81ff0681",
   390 => x"16585473",
   391 => x"802e8a38",
   392 => x"9c5380c3",
   393 => x"c4528caf",
   394 => x"048b53bc",
   395 => x"8c0852bc",
   396 => x"be16518c",
   397 => x"e6047416",
   398 => x"822b8ac2",
   399 => x"0bba8c12",
   400 => x"0c547681",
   401 => x"ff068116",
   402 => x"58547380",
   403 => x"2e8a389c",
   404 => x"5380c3c4",
   405 => x"528cde04",
   406 => x"8b53bc8c",
   407 => x"08527775",
   408 => x"3110bcbc",
   409 => x"05517655",
   410 => x"89cf2d8c",
   411 => x"ff047490",
   412 => x"29753170",
   413 => x"10bcbc05",
   414 => x"5154bc8c",
   415 => x"08743481",
   416 => x"1959748b",
   417 => x"24a0388b",
   418 => x"bd047490",
   419 => x"29753170",
   420 => x"10bcbc05",
   421 => x"8c773157",
   422 => x"51548074",
   423 => x"349e14ff",
   424 => x"16565474",
   425 => x"f53802a4",
   426 => x"050d0402",
   427 => x"fc050dbb",
   428 => x"b8081351",
   429 => x"89f82dbc",
   430 => x"8c08802e",
   431 => x"8838bc8c",
   432 => x"08519281",
   433 => x"2d800bbb",
   434 => x"b80c8afc",
   435 => x"2dab9e2d",
   436 => x"0284050d",
   437 => x"0402fc05",
   438 => x"0d725170",
   439 => x"fd2ead38",
   440 => x"70fd248a",
   441 => x"3870fc2e",
   442 => x"80c4388e",
   443 => x"b60470fe",
   444 => x"2eb13870",
   445 => x"ff2e0981",
   446 => x"06bc38bb",
   447 => x"b8085170",
   448 => x"802eb338",
   449 => x"ff11bbb8",
   450 => x"0c8eb604",
   451 => x"bbb808f0",
   452 => x"0570bbb8",
   453 => x"0c517080",
   454 => x"259c3880",
   455 => x"0bbbb80c",
   456 => x"8eb604bb",
   457 => x"b8088105",
   458 => x"bbb80c8e",
   459 => x"b604bbb8",
   460 => x"089005bb",
   461 => x"b80c8afc",
   462 => x"2dab9e2d",
   463 => x"0284050d",
   464 => x"0402fc05",
   465 => x"0dbcb408",
   466 => x"fb06bcb4",
   467 => x"0c72518a",
   468 => x"c22d0284",
   469 => x"050d0402",
   470 => x"fc050dbc",
   471 => x"b4088407",
   472 => x"bcb40c72",
   473 => x"518ac22d",
   474 => x"0284050d",
   475 => x"0402fc05",
   476 => x"0d800bbb",
   477 => x"b80c8afc",
   478 => x"2dba8451",
   479 => x"acbd2db9",
   480 => x"ec51acd0",
   481 => x"2d028405",
   482 => x"0d0402f8",
   483 => x"050d80c6",
   484 => x"b0088206",
   485 => x"b99c3352",
   486 => x"5270802e",
   487 => x"85387181",
   488 => x"0752b9b4",
   489 => x"33517080",
   490 => x"2e853871",
   491 => x"840752bc",
   492 => x"b808802e",
   493 => x"85387190",
   494 => x"075271bc",
   495 => x"8c0c0288",
   496 => x"050d0402",
   497 => x"f4050d81",
   498 => x"0bbcb80c",
   499 => x"90518694",
   500 => x"2d810bfe",
   501 => x"c40c900b",
   502 => x"fec00c84",
   503 => x"0bfec40c",
   504 => x"830bfecc",
   505 => x"0ca8aa2d",
   506 => x"aac02da8",
   507 => x"8d2da88d",
   508 => x"2d81fb2d",
   509 => x"815184e9",
   510 => x"2da88d2d",
   511 => x"a88d2d81",
   512 => x"5184e92d",
   513 => x"0b0b0bb7",
   514 => x"9c5185f5",
   515 => x"2d8452a2",
   516 => x"9a2d939e",
   517 => x"2dbc8c08",
   518 => x"802e8638",
   519 => x"fe5290a9",
   520 => x"04ff1252",
   521 => x"718024e7",
   522 => x"3871802e",
   523 => x"81863886",
   524 => x"c12d0b0b",
   525 => x"0bb7b451",
   526 => x"87be2dbc",
   527 => x"8c08802e",
   528 => x"8f38b8fc",
   529 => x"51acbd2d",
   530 => x"805184e9",
   531 => x"2d90da04",
   532 => x"bc8c0851",
   533 => x"8eed2daa",
   534 => x"cc2da8c3",
   535 => x"2dacd62d",
   536 => x"bc8c0880",
   537 => x"c6b40888",
   538 => x"2b80c6b8",
   539 => x"0807fed8",
   540 => x"0c538f8a",
   541 => x"2dbc8c08",
   542 => x"bcb4082e",
   543 => x"a238bc8c",
   544 => x"08bcb40c",
   545 => x"bc8c08fe",
   546 => x"c00c8452",
   547 => x"725184e9",
   548 => x"2da88d2d",
   549 => x"a88d2dff",
   550 => x"12527180",
   551 => x"25ee3872",
   552 => x"802e8938",
   553 => x"8a0bfec4",
   554 => x"0c90da04",
   555 => x"820bfec4",
   556 => x"0c90da04",
   557 => x"0b0b0bb7",
   558 => x"c05185f5",
   559 => x"2d800bbc",
   560 => x"8c0c028c",
   561 => x"050d0402",
   562 => x"e8050d77",
   563 => x"797b5855",
   564 => x"55805372",
   565 => x"76259f38",
   566 => x"74708105",
   567 => x"56337470",
   568 => x"81055633",
   569 => x"52527171",
   570 => x"2e863881",
   571 => x"5191f804",
   572 => x"81135391",
   573 => x"d3048051",
   574 => x"70bc8c0c",
   575 => x"0298050d",
   576 => x"0402ec05",
   577 => x"0d765574",
   578 => x"802eba38",
   579 => x"9a152251",
   580 => x"a6d42dbc",
   581 => x"8c08bc8c",
   582 => x"0880c5f4",
   583 => x"0cbc8c08",
   584 => x"545480c5",
   585 => x"d008802e",
   586 => x"97389415",
   587 => x"2251a6d4",
   588 => x"2dbc8c08",
   589 => x"902b83ff",
   590 => x"f00a0670",
   591 => x"75075153",
   592 => x"7280c5f4",
   593 => x"0c80c5f4",
   594 => x"08537280",
   595 => x"2e9d3880",
   596 => x"c5c808fe",
   597 => x"14712980",
   598 => x"c5dc0805",
   599 => x"80c5f80c",
   600 => x"70842b80",
   601 => x"c5d40c54",
   602 => x"93990480",
   603 => x"c5e00880",
   604 => x"c5f40c80",
   605 => x"c5e40880",
   606 => x"c5f80c80",
   607 => x"c5d00880",
   608 => x"2e8b3880",
   609 => x"c5c80884",
   610 => x"2b539394",
   611 => x"0480c5e8",
   612 => x"08842b53",
   613 => x"7280c5d4",
   614 => x"0c029405",
   615 => x"0d0402d8",
   616 => x"050d800b",
   617 => x"80c5d00c",
   618 => x"bfc45280",
   619 => x"51a5842d",
   620 => x"bc8c0854",
   621 => x"bc8c088c",
   622 => x"38b7d451",
   623 => x"85f52d73",
   624 => x"55989104",
   625 => x"8056810b",
   626 => x"80c5fc0c",
   627 => x"8853b7e0",
   628 => x"52bffa51",
   629 => x"91c72dbc",
   630 => x"8c08762e",
   631 => x"09810688",
   632 => x"38bc8c08",
   633 => x"80c5fc0c",
   634 => x"8853b7ec",
   635 => x"5280c096",
   636 => x"5191c72d",
   637 => x"bc8c0888",
   638 => x"38bc8c08",
   639 => x"80c5fc0c",
   640 => x"80c5fc08",
   641 => x"802e80ea",
   642 => x"3880c38a",
   643 => x"3380c38b",
   644 => x"3371982b",
   645 => x"71902b07",
   646 => x"80c38c33",
   647 => x"70882b72",
   648 => x"0780c38d",
   649 => x"33710780",
   650 => x"c3c23380",
   651 => x"c3c33371",
   652 => x"882b0753",
   653 => x"5f54525a",
   654 => x"56575573",
   655 => x"81abaa2e",
   656 => x"0981068d",
   657 => x"387551a6",
   658 => x"a42dbc8c",
   659 => x"085694de",
   660 => x"047382d4",
   661 => x"d52e8738",
   662 => x"b7f85195",
   663 => x"a104bfc4",
   664 => x"527551a5",
   665 => x"842dbc8c",
   666 => x"0855bc8c",
   667 => x"08802e83",
   668 => x"a0388853",
   669 => x"b7ec5280",
   670 => x"c0965191",
   671 => x"c72dbc8c",
   672 => x"088a3881",
   673 => x"0b80c5d0",
   674 => x"0c95a704",
   675 => x"8853b7e0",
   676 => x"52bffa51",
   677 => x"91c72dbc",
   678 => x"8c08802e",
   679 => x"8a38b88c",
   680 => x"5185f52d",
   681 => x"95f30480",
   682 => x"c3c23354",
   683 => x"7380d52e",
   684 => x"098106bf",
   685 => x"3880c3c3",
   686 => x"33547381",
   687 => x"aa2e0981",
   688 => x"06b13880",
   689 => x"0bbfc433",
   690 => x"56547481",
   691 => x"e92e8338",
   692 => x"81547481",
   693 => x"eb2e8c38",
   694 => x"80557375",
   695 => x"2e098106",
   696 => x"82af38bf",
   697 => x"cf335574",
   698 => x"8a38bfd0",
   699 => x"33547382",
   700 => x"2e863880",
   701 => x"55989104",
   702 => x"bfd13370",
   703 => x"80c5c80c",
   704 => x"ff0580c5",
   705 => x"cc0cbfd2",
   706 => x"33bfd333",
   707 => x"58760577",
   708 => x"82802905",
   709 => x"7080c5d8",
   710 => x"0cbfd433",
   711 => x"7080c5ec",
   712 => x"0c80c5d0",
   713 => x"08595758",
   714 => x"76802e81",
   715 => x"95388853",
   716 => x"b7ec5280",
   717 => x"c0965191",
   718 => x"c72dbc8c",
   719 => x"0881d238",
   720 => x"80c5c808",
   721 => x"70842b80",
   722 => x"c5d40c70",
   723 => x"80c5e80c",
   724 => x"bfe933bf",
   725 => x"e8337182",
   726 => x"802905bf",
   727 => x"ea337084",
   728 => x"80802912",
   729 => x"bfeb3370",
   730 => x"81800a29",
   731 => x"127080c5",
   732 => x"f00c80c5",
   733 => x"ec087129",
   734 => x"80c5d808",
   735 => x"057080c5",
   736 => x"dc0cbff1",
   737 => x"33bff033",
   738 => x"71828029",
   739 => x"05bff233",
   740 => x"70848080",
   741 => x"2912bff3",
   742 => x"3370982b",
   743 => x"81f00a06",
   744 => x"72057080",
   745 => x"c5e00cfe",
   746 => x"117e2977",
   747 => x"0580c5e4",
   748 => x"0c525952",
   749 => x"43545e51",
   750 => x"5259525d",
   751 => x"57595798",
   752 => x"8a04bfd6",
   753 => x"33bfd533",
   754 => x"71828029",
   755 => x"057080c5",
   756 => x"d40c70a0",
   757 => x"2983ff05",
   758 => x"70892a70",
   759 => x"80c5e80c",
   760 => x"bfdb33bf",
   761 => x"da337182",
   762 => x"80290570",
   763 => x"80c5f00c",
   764 => x"7b71291e",
   765 => x"7080c5e4",
   766 => x"0c7d80c5",
   767 => x"e00c7305",
   768 => x"80c5dc0c",
   769 => x"555e5151",
   770 => x"55558051",
   771 => x"92812d81",
   772 => x"5574bc8c",
   773 => x"0c02a805",
   774 => x"0d0402ec",
   775 => x"050d7670",
   776 => x"872c7180",
   777 => x"ff065556",
   778 => x"5480c5d0",
   779 => x"088a3873",
   780 => x"882c7481",
   781 => x"ff065455",
   782 => x"bfc45280",
   783 => x"c5d80815",
   784 => x"51a5842d",
   785 => x"bc8c0854",
   786 => x"bc8c0880",
   787 => x"2eb23880",
   788 => x"c5d00880",
   789 => x"2e983872",
   790 => x"8429bfc4",
   791 => x"05700852",
   792 => x"53a6a42d",
   793 => x"bc8c08f0",
   794 => x"0a065398",
   795 => x"fe047210",
   796 => x"bfc40570",
   797 => x"225253a6",
   798 => x"d42dbc8c",
   799 => x"08537254",
   800 => x"73bc8c0c",
   801 => x"0294050d",
   802 => x"0402e005",
   803 => x"0d797084",
   804 => x"2c80c5f8",
   805 => x"0805718f",
   806 => x"06525553",
   807 => x"728938bf",
   808 => x"c4527351",
   809 => x"a5842d72",
   810 => x"a029bfc4",
   811 => x"05548074",
   812 => x"33565374",
   813 => x"732e8338",
   814 => x"81537481",
   815 => x"e52e81b8",
   816 => x"38817074",
   817 => x"06545872",
   818 => x"802e81ac",
   819 => x"388b1433",
   820 => x"70832a79",
   821 => x"06585676",
   822 => x"9638bbbc",
   823 => x"08537286",
   824 => x"387280c3",
   825 => x"c43476bb",
   826 => x"bc0c7353",
   827 => x"9afa0475",
   828 => x"8f2e0981",
   829 => x"06818138",
   830 => x"749f068d",
   831 => x"2980c3b7",
   832 => x"11515381",
   833 => x"14337370",
   834 => x"81055534",
   835 => x"83143373",
   836 => x"70810555",
   837 => x"34851433",
   838 => x"73708105",
   839 => x"55348714",
   840 => x"33737081",
   841 => x"05553489",
   842 => x"14337370",
   843 => x"81055534",
   844 => x"8e143373",
   845 => x"70810555",
   846 => x"34901433",
   847 => x"73708105",
   848 => x"55349214",
   849 => x"33737081",
   850 => x"05553494",
   851 => x"14337370",
   852 => x"81055534",
   853 => x"96143373",
   854 => x"70810555",
   855 => x"34981433",
   856 => x"73708105",
   857 => x"55349c14",
   858 => x"33737081",
   859 => x"0555349e",
   860 => x"14337334",
   861 => x"77bbbc0c",
   862 => x"805372bc",
   863 => x"8c0c02a0",
   864 => x"050d0402",
   865 => x"cc050d7e",
   866 => x"605e5a80",
   867 => x"0b80c5f4",
   868 => x"0880c5f8",
   869 => x"08595c56",
   870 => x"805880c5",
   871 => x"d408782e",
   872 => x"81a83877",
   873 => x"8f06a017",
   874 => x"5754738f",
   875 => x"38bfc452",
   876 => x"76518117",
   877 => x"57a5842d",
   878 => x"bfc45680",
   879 => x"76335654",
   880 => x"74742e83",
   881 => x"38815474",
   882 => x"81e52e80",
   883 => x"f1388170",
   884 => x"7506555c",
   885 => x"73802e80",
   886 => x"e5388b16",
   887 => x"33980659",
   888 => x"7880db38",
   889 => x"8b537c52",
   890 => x"755191c7",
   891 => x"2dbc8c08",
   892 => x"80cc389c",
   893 => x"160851a6",
   894 => x"a42dbc8c",
   895 => x"08841b0c",
   896 => x"9a162251",
   897 => x"a6d42dbc",
   898 => x"8c08bc8c",
   899 => x"08881c0c",
   900 => x"bc8c0855",
   901 => x"5580c5d0",
   902 => x"08802e96",
   903 => x"38941622",
   904 => x"51a6d42d",
   905 => x"bc8c0890",
   906 => x"2b83fff0",
   907 => x"0a067016",
   908 => x"51547388",
   909 => x"1b0c787a",
   910 => x"0c7b549d",
   911 => x"83048118",
   912 => x"5880c5d4",
   913 => x"087826fe",
   914 => x"da3880c5",
   915 => x"d008802e",
   916 => x"b0387a51",
   917 => x"989a2dbc",
   918 => x"8c08bc8c",
   919 => x"0880ffff",
   920 => x"fff80655",
   921 => x"5b7380ff",
   922 => x"fffff82e",
   923 => x"9438bc8c",
   924 => x"08fe0580",
   925 => x"c5c80829",
   926 => x"80c5dc08",
   927 => x"05579b98",
   928 => x"04805473",
   929 => x"bc8c0c02",
   930 => x"b4050d04",
   931 => x"02f4050d",
   932 => x"74700881",
   933 => x"05710c70",
   934 => x"0880c5cc",
   935 => x"08065353",
   936 => x"718e3888",
   937 => x"13085198",
   938 => x"9a2dbc8c",
   939 => x"0888140c",
   940 => x"810bbc8c",
   941 => x"0c028c05",
   942 => x"0d0402f0",
   943 => x"050d7588",
   944 => x"1108fe05",
   945 => x"80c5c808",
   946 => x"2980c5dc",
   947 => x"08117208",
   948 => x"80c5cc08",
   949 => x"06057955",
   950 => x"535454a5",
   951 => x"842d0290",
   952 => x"050d0402",
   953 => x"f0050d75",
   954 => x"881108fe",
   955 => x"0580c5c8",
   956 => x"082980c5",
   957 => x"dc081172",
   958 => x"0880c5cc",
   959 => x"08060579",
   960 => x"55535454",
   961 => x"a3c42d02",
   962 => x"90050d04",
   963 => x"02f4050d",
   964 => x"d45281ff",
   965 => x"720c7108",
   966 => x"5381ff72",
   967 => x"0c72882b",
   968 => x"83fe8006",
   969 => x"72087081",
   970 => x"ff065152",
   971 => x"5381ff72",
   972 => x"0c727107",
   973 => x"882b7208",
   974 => x"7081ff06",
   975 => x"51525381",
   976 => x"ff720c72",
   977 => x"7107882b",
   978 => x"72087081",
   979 => x"ff067207",
   980 => x"bc8c0c52",
   981 => x"53028c05",
   982 => x"0d0402f4",
   983 => x"050d7476",
   984 => x"7181ff06",
   985 => x"d40c5353",
   986 => x"80c68008",
   987 => x"85387189",
   988 => x"2b527198",
   989 => x"2ad40c71",
   990 => x"902a7081",
   991 => x"ff06d40c",
   992 => x"5171882a",
   993 => x"7081ff06",
   994 => x"d40c5171",
   995 => x"81ff06d4",
   996 => x"0c72902a",
   997 => x"7081ff06",
   998 => x"d40c51d4",
   999 => x"087081ff",
  1000 => x"06515182",
  1001 => x"b8bf5270",
  1002 => x"81ff2e09",
  1003 => x"81069438",
  1004 => x"81ff0bd4",
  1005 => x"0cd40870",
  1006 => x"81ff06ff",
  1007 => x"14545151",
  1008 => x"71e53870",
  1009 => x"bc8c0c02",
  1010 => x"8c050d04",
  1011 => x"02fc050d",
  1012 => x"81c75181",
  1013 => x"ff0bd40c",
  1014 => x"ff115170",
  1015 => x"8025f438",
  1016 => x"0284050d",
  1017 => x"0402f005",
  1018 => x"0d9fcc2d",
  1019 => x"8fcf5380",
  1020 => x"5287fc80",
  1021 => x"f7519eda",
  1022 => x"2dbc8c08",
  1023 => x"54bc8c08",
  1024 => x"812e0981",
  1025 => x"06a33881",
  1026 => x"ff0bd40c",
  1027 => x"820a5284",
  1028 => x"9c80e951",
  1029 => x"9eda2dbc",
  1030 => x"8c088b38",
  1031 => x"81ff0bd4",
  1032 => x"0c7353a0",
  1033 => x"af049fcc",
  1034 => x"2dff1353",
  1035 => x"72c13872",
  1036 => x"bc8c0c02",
  1037 => x"90050d04",
  1038 => x"02f4050d",
  1039 => x"81ff0bd4",
  1040 => x"0c935380",
  1041 => x"5287fc80",
  1042 => x"c1519eda",
  1043 => x"2dbc8c08",
  1044 => x"8b3881ff",
  1045 => x"0bd40c81",
  1046 => x"53a0e504",
  1047 => x"9fcc2dff",
  1048 => x"135372df",
  1049 => x"3872bc8c",
  1050 => x"0c028c05",
  1051 => x"0d0402f0",
  1052 => x"050d9fcc",
  1053 => x"2d83aa52",
  1054 => x"849c80c8",
  1055 => x"519eda2d",
  1056 => x"bc8c0881",
  1057 => x"2e098106",
  1058 => x"92389e8c",
  1059 => x"2dbc8c08",
  1060 => x"83ffff06",
  1061 => x"537283aa",
  1062 => x"2e9738a0",
  1063 => x"b82da1ac",
  1064 => x"048154a2",
  1065 => x"9104b898",
  1066 => x"5185f52d",
  1067 => x"8054a291",
  1068 => x"0481ff0b",
  1069 => x"d40cb153",
  1070 => x"9fe52dbc",
  1071 => x"8c08802e",
  1072 => x"80c03880",
  1073 => x"5287fc80",
  1074 => x"fa519eda",
  1075 => x"2dbc8c08",
  1076 => x"b13881ff",
  1077 => x"0bd40cd4",
  1078 => x"085381ff",
  1079 => x"0bd40c81",
  1080 => x"ff0bd40c",
  1081 => x"81ff0bd4",
  1082 => x"0c81ff0b",
  1083 => x"d40c7286",
  1084 => x"2a708106",
  1085 => x"bc8c0856",
  1086 => x"51537280",
  1087 => x"2e9338a1",
  1088 => x"a1047282",
  1089 => x"2eff9f38",
  1090 => x"ff135372",
  1091 => x"ffaa3872",
  1092 => x"5473bc8c",
  1093 => x"0c029005",
  1094 => x"0d0402f0",
  1095 => x"050d810b",
  1096 => x"80c6800c",
  1097 => x"8454d008",
  1098 => x"708f2a70",
  1099 => x"81065151",
  1100 => x"5372f338",
  1101 => x"72d00c9f",
  1102 => x"cc2db8a8",
  1103 => x"5185f52d",
  1104 => x"d008708f",
  1105 => x"2a708106",
  1106 => x"51515372",
  1107 => x"f338810b",
  1108 => x"d00cb153",
  1109 => x"805284d4",
  1110 => x"80c0519e",
  1111 => x"da2dbc8c",
  1112 => x"08812ea1",
  1113 => x"3872822e",
  1114 => x"0981068c",
  1115 => x"38b8b451",
  1116 => x"85f52d80",
  1117 => x"53a3bb04",
  1118 => x"ff135372",
  1119 => x"d738ff14",
  1120 => x"5473ffa2",
  1121 => x"38a0ee2d",
  1122 => x"bc8c0880",
  1123 => x"c6800cbc",
  1124 => x"8c088b38",
  1125 => x"815287fc",
  1126 => x"80d0519e",
  1127 => x"da2d81ff",
  1128 => x"0bd40cd0",
  1129 => x"08708f2a",
  1130 => x"70810651",
  1131 => x"515372f3",
  1132 => x"3872d00c",
  1133 => x"81ff0bd4",
  1134 => x"0c815372",
  1135 => x"bc8c0c02",
  1136 => x"90050d04",
  1137 => x"02e8050d",
  1138 => x"785681ff",
  1139 => x"0bd40cd0",
  1140 => x"08708f2a",
  1141 => x"70810651",
  1142 => x"515372f3",
  1143 => x"3882810b",
  1144 => x"d00c81ff",
  1145 => x"0bd40c77",
  1146 => x"5287fc80",
  1147 => x"d8519eda",
  1148 => x"2dbc8c08",
  1149 => x"802e8c38",
  1150 => x"b8cc5185",
  1151 => x"f52d8153",
  1152 => x"a4fb0481",
  1153 => x"ff0bd40c",
  1154 => x"81fe0bd4",
  1155 => x"0c80ff55",
  1156 => x"75708405",
  1157 => x"57087098",
  1158 => x"2ad40c70",
  1159 => x"902c7081",
  1160 => x"ff06d40c",
  1161 => x"5470882c",
  1162 => x"7081ff06",
  1163 => x"d40c5470",
  1164 => x"81ff06d4",
  1165 => x"0c54ff15",
  1166 => x"55748025",
  1167 => x"d33881ff",
  1168 => x"0bd40c81",
  1169 => x"ff0bd40c",
  1170 => x"81ff0bd4",
  1171 => x"0c868da0",
  1172 => x"5481ff0b",
  1173 => x"d40cd408",
  1174 => x"81ff0655",
  1175 => x"748738ff",
  1176 => x"145473ed",
  1177 => x"3881ff0b",
  1178 => x"d40cd008",
  1179 => x"708f2a70",
  1180 => x"81065151",
  1181 => x"5372f338",
  1182 => x"72d00c72",
  1183 => x"bc8c0c02",
  1184 => x"98050d04",
  1185 => x"02e8050d",
  1186 => x"78558056",
  1187 => x"81ff0bd4",
  1188 => x"0cd00870",
  1189 => x"8f2a7081",
  1190 => x"06515153",
  1191 => x"72f33882",
  1192 => x"810bd00c",
  1193 => x"81ff0bd4",
  1194 => x"0c775287",
  1195 => x"fc80d151",
  1196 => x"9eda2d80",
  1197 => x"dbc6df54",
  1198 => x"bc8c0880",
  1199 => x"2e8a38b8",
  1200 => x"dc5185f5",
  1201 => x"2da69b04",
  1202 => x"81ff0bd4",
  1203 => x"0cd40870",
  1204 => x"81ff0651",
  1205 => x"537281fe",
  1206 => x"2e098106",
  1207 => x"9d3880ff",
  1208 => x"539e8c2d",
  1209 => x"bc8c0875",
  1210 => x"70840557",
  1211 => x"0cff1353",
  1212 => x"728025ed",
  1213 => x"388156a6",
  1214 => x"8004ff14",
  1215 => x"5473c938",
  1216 => x"81ff0bd4",
  1217 => x"0c81ff0b",
  1218 => x"d40cd008",
  1219 => x"708f2a70",
  1220 => x"81065151",
  1221 => x"5372f338",
  1222 => x"72d00c75",
  1223 => x"bc8c0c02",
  1224 => x"98050d04",
  1225 => x"02f4050d",
  1226 => x"7470882a",
  1227 => x"83fe8006",
  1228 => x"7072982a",
  1229 => x"0772882b",
  1230 => x"87fc8080",
  1231 => x"0673982b",
  1232 => x"81f00a06",
  1233 => x"71730707",
  1234 => x"bc8c0c56",
  1235 => x"51535102",
  1236 => x"8c050d04",
  1237 => x"02f8050d",
  1238 => x"028e0533",
  1239 => x"74882b07",
  1240 => x"7083ffff",
  1241 => x"06bc8c0c",
  1242 => x"51028805",
  1243 => x"0d0402fc",
  1244 => x"050d7251",
  1245 => x"80710c80",
  1246 => x"0b84120c",
  1247 => x"0284050d",
  1248 => x"0402f005",
  1249 => x"0d757008",
  1250 => x"84120853",
  1251 => x"5353ff54",
  1252 => x"71712ea8",
  1253 => x"38aac62d",
  1254 => x"84130870",
  1255 => x"84291488",
  1256 => x"11700870",
  1257 => x"81ff0684",
  1258 => x"18088111",
  1259 => x"8706841a",
  1260 => x"0c535155",
  1261 => x"515151aa",
  1262 => x"c02d7154",
  1263 => x"73bc8c0c",
  1264 => x"0290050d",
  1265 => x"0402f805",
  1266 => x"0daac62d",
  1267 => x"e008708b",
  1268 => x"2a708106",
  1269 => x"51525270",
  1270 => x"802ea138",
  1271 => x"80c68408",
  1272 => x"70842980",
  1273 => x"c68c0573",
  1274 => x"81ff0671",
  1275 => x"0c515180",
  1276 => x"c6840881",
  1277 => x"11870680",
  1278 => x"c6840c51",
  1279 => x"800b80c6",
  1280 => x"ac0caab9",
  1281 => x"2daac02d",
  1282 => x"0288050d",
  1283 => x"0402fc05",
  1284 => x"0daac62d",
  1285 => x"810b80c6",
  1286 => x"ac0caac0",
  1287 => x"2d80c6ac",
  1288 => x"085170f9",
  1289 => x"38028405",
  1290 => x"0d0402fc",
  1291 => x"050d80c6",
  1292 => x"8451a6ee",
  1293 => x"2da7c551",
  1294 => x"aab42da9",
  1295 => x"de2d0284",
  1296 => x"050d0402",
  1297 => x"f4050da9",
  1298 => x"c504bc8c",
  1299 => x"0881f02e",
  1300 => x"09810689",
  1301 => x"38810bbc",
  1302 => x"800ca9c5",
  1303 => x"04bc8c08",
  1304 => x"81e02e09",
  1305 => x"81068938",
  1306 => x"810bbc84",
  1307 => x"0ca9c504",
  1308 => x"bc8c0852",
  1309 => x"bc840880",
  1310 => x"2e8838bc",
  1311 => x"8c088180",
  1312 => x"05527184",
  1313 => x"2c728f06",
  1314 => x"5353bc80",
  1315 => x"08802e99",
  1316 => x"38728429",
  1317 => x"bbc00572",
  1318 => x"1381712b",
  1319 => x"70097308",
  1320 => x"06730c51",
  1321 => x"5353a9bb",
  1322 => x"04728429",
  1323 => x"bbc00572",
  1324 => x"1383712b",
  1325 => x"72080772",
  1326 => x"0c535380",
  1327 => x"0bbc840c",
  1328 => x"800bbc80",
  1329 => x"0c80c684",
  1330 => x"51a7812d",
  1331 => x"bc8c08ff",
  1332 => x"24fef738",
  1333 => x"800bbc8c",
  1334 => x"0c028c05",
  1335 => x"0d0402f8",
  1336 => x"050dbbc0",
  1337 => x"528f5180",
  1338 => x"72708405",
  1339 => x"540cff11",
  1340 => x"51708025",
  1341 => x"f2380288",
  1342 => x"050d0402",
  1343 => x"f0050d75",
  1344 => x"51aac62d",
  1345 => x"70822cfc",
  1346 => x"06bbc011",
  1347 => x"72109e06",
  1348 => x"71087072",
  1349 => x"2a708306",
  1350 => x"82742b70",
  1351 => x"09740676",
  1352 => x"0c545156",
  1353 => x"57535153",
  1354 => x"aac02d71",
  1355 => x"bc8c0c02",
  1356 => x"90050d04",
  1357 => x"7180cc0c",
  1358 => x"04ffb008",
  1359 => x"bc8c0c04",
  1360 => x"810bffb0",
  1361 => x"0c04800b",
  1362 => x"ffb00c04",
  1363 => x"02fc050d",
  1364 => x"810bbc88",
  1365 => x"0c815184",
  1366 => x"e92d0284",
  1367 => x"050d0402",
  1368 => x"fc050d80",
  1369 => x"0bbc880c",
  1370 => x"805184e9",
  1371 => x"2d028405",
  1372 => x"0d0402ec",
  1373 => x"050d7654",
  1374 => x"8052870b",
  1375 => x"88153356",
  1376 => x"53747224",
  1377 => x"8338a053",
  1378 => x"725182f2",
  1379 => x"2d81128b",
  1380 => x"15335452",
  1381 => x"727225e2",
  1382 => x"38029405",
  1383 => x"0d0402f0",
  1384 => x"050d80c6",
  1385 => x"bc085481",
  1386 => x"fb2d800b",
  1387 => x"80c6c00c",
  1388 => x"7308802e",
  1389 => x"81823882",
  1390 => x"0bbca00c",
  1391 => x"80c6c008",
  1392 => x"8f06bc9c",
  1393 => x"0c730852",
  1394 => x"71832e96",
  1395 => x"38718326",
  1396 => x"89387181",
  1397 => x"2ead38ac",
  1398 => x"a1047185",
  1399 => x"2e9d38ac",
  1400 => x"a1048814",
  1401 => x"33841508",
  1402 => x"b8ec5354",
  1403 => x"5285f52d",
  1404 => x"71842913",
  1405 => x"70085252",
  1406 => x"aca50473",
  1407 => x"51aaf22d",
  1408 => x"aca10480",
  1409 => x"c6b00888",
  1410 => x"15082c70",
  1411 => x"81065152",
  1412 => x"71802e87",
  1413 => x"38b8f051",
  1414 => x"ac9e04b8",
  1415 => x"f45185f5",
  1416 => x"2d841408",
  1417 => x"5185f52d",
  1418 => x"80c6c008",
  1419 => x"810580c6",
  1420 => x"c00c8c14",
  1421 => x"54abb004",
  1422 => x"0290050d",
  1423 => x"047180c6",
  1424 => x"bc0cab9e",
  1425 => x"2d80c6c0",
  1426 => x"08ff0580",
  1427 => x"c6c40c04",
  1428 => x"7180c6c8",
  1429 => x"0c0402e8",
  1430 => x"050d80c6",
  1431 => x"bc0880c6",
  1432 => x"c8085755",
  1433 => x"80f851a9",
  1434 => x"fb2dbc8c",
  1435 => x"08812a70",
  1436 => x"81065152",
  1437 => x"719b3887",
  1438 => x"51a9fb2d",
  1439 => x"bc8c0881",
  1440 => x"2a708106",
  1441 => x"51527180",
  1442 => x"2eb138ad",
  1443 => x"9104a8c3",
  1444 => x"2d8751a9",
  1445 => x"fb2dbc8c",
  1446 => x"08f438ad",
  1447 => x"a104a8c3",
  1448 => x"2d80f851",
  1449 => x"a9fb2dbc",
  1450 => x"8c08f338",
  1451 => x"bc880881",
  1452 => x"3270bc88",
  1453 => x"0c705252",
  1454 => x"84e92d80",
  1455 => x"0b80c6b4",
  1456 => x"0c800b80",
  1457 => x"c6b80cbc",
  1458 => x"880882fd",
  1459 => x"3880da51",
  1460 => x"a9fb2dbc",
  1461 => x"8c08802e",
  1462 => x"8c3880c6",
  1463 => x"b4088180",
  1464 => x"0780c6b4",
  1465 => x"0c80d951",
  1466 => x"a9fb2dbc",
  1467 => x"8c08802e",
  1468 => x"8c3880c6",
  1469 => x"b40880c0",
  1470 => x"0780c6b4",
  1471 => x"0c819451",
  1472 => x"a9fb2dbc",
  1473 => x"8c08802e",
  1474 => x"8b3880c6",
  1475 => x"b4089007",
  1476 => x"80c6b40c",
  1477 => x"819151a9",
  1478 => x"fb2dbc8c",
  1479 => x"08802e8b",
  1480 => x"3880c6b4",
  1481 => x"08a00780",
  1482 => x"c6b40c81",
  1483 => x"f551a9fb",
  1484 => x"2dbc8c08",
  1485 => x"802e8b38",
  1486 => x"80c6b408",
  1487 => x"810780c6",
  1488 => x"b40c81f2",
  1489 => x"51a9fb2d",
  1490 => x"bc8c0880",
  1491 => x"2e8b3880",
  1492 => x"c6b40882",
  1493 => x"0780c6b4",
  1494 => x"0c81eb51",
  1495 => x"a9fb2dbc",
  1496 => x"8c08802e",
  1497 => x"8b3880c6",
  1498 => x"b4088407",
  1499 => x"80c6b40c",
  1500 => x"81f451a9",
  1501 => x"fb2dbc8c",
  1502 => x"08802e8b",
  1503 => x"3880c6b4",
  1504 => x"08880780",
  1505 => x"c6b40c80",
  1506 => x"d851a9fb",
  1507 => x"2dbc8c08",
  1508 => x"802e8c38",
  1509 => x"80c6b808",
  1510 => x"81800780",
  1511 => x"c6b80c92",
  1512 => x"51a9fb2d",
  1513 => x"bc8c0880",
  1514 => x"2e8c3880",
  1515 => x"c6b80880",
  1516 => x"c00780c6",
  1517 => x"b80c9451",
  1518 => x"a9fb2dbc",
  1519 => x"8c08802e",
  1520 => x"8b3880c6",
  1521 => x"b8089007",
  1522 => x"80c6b80c",
  1523 => x"9151a9fb",
  1524 => x"2dbc8c08",
  1525 => x"802e8b38",
  1526 => x"80c6b808",
  1527 => x"a00780c6",
  1528 => x"b80c9d51",
  1529 => x"a9fb2dbc",
  1530 => x"8c08802e",
  1531 => x"8b3880c6",
  1532 => x"b8088107",
  1533 => x"80c6b80c",
  1534 => x"9b51a9fb",
  1535 => x"2dbc8c08",
  1536 => x"802e8b38",
  1537 => x"80c6b808",
  1538 => x"820780c6",
  1539 => x"b80c9c51",
  1540 => x"a9fb2dbc",
  1541 => x"8c08802e",
  1542 => x"8b3880c6",
  1543 => x"b8088407",
  1544 => x"80c6b80c",
  1545 => x"a351a9fb",
  1546 => x"2dbc8c08",
  1547 => x"802e8b38",
  1548 => x"80c6b808",
  1549 => x"880780c6",
  1550 => x"b80c81fd",
  1551 => x"51a9fb2d",
  1552 => x"81fa51a9",
  1553 => x"fb2db5fd",
  1554 => x"0481f551",
  1555 => x"a9fb2dbc",
  1556 => x"8c08812a",
  1557 => x"70810651",
  1558 => x"5271802e",
  1559 => x"b33880c6",
  1560 => x"c4085271",
  1561 => x"802e8a38",
  1562 => x"ff1280c6",
  1563 => x"c40cb190",
  1564 => x"0480c6c0",
  1565 => x"081080c6",
  1566 => x"c0080570",
  1567 => x"84291651",
  1568 => x"52881208",
  1569 => x"802e8938",
  1570 => x"ff518812",
  1571 => x"0852712d",
  1572 => x"81f251a9",
  1573 => x"fb2dbc8c",
  1574 => x"08812a70",
  1575 => x"81065152",
  1576 => x"71802eb4",
  1577 => x"3880c6c0",
  1578 => x"08ff1180",
  1579 => x"c6c40856",
  1580 => x"53537372",
  1581 => x"258a3881",
  1582 => x"1480c6c4",
  1583 => x"0cb1d804",
  1584 => x"72101370",
  1585 => x"84291651",
  1586 => x"52881208",
  1587 => x"802e8938",
  1588 => x"fe518812",
  1589 => x"0852712d",
  1590 => x"81fd51a9",
  1591 => x"fb2dbc8c",
  1592 => x"08812a70",
  1593 => x"81065152",
  1594 => x"71802eb1",
  1595 => x"3880c6c4",
  1596 => x"08802e8a",
  1597 => x"38800b80",
  1598 => x"c6c40cb2",
  1599 => x"9d0480c6",
  1600 => x"c0081080",
  1601 => x"c6c00805",
  1602 => x"70842916",
  1603 => x"51528812",
  1604 => x"08802e89",
  1605 => x"38fd5188",
  1606 => x"12085271",
  1607 => x"2d81fa51",
  1608 => x"a9fb2dbc",
  1609 => x"8c08812a",
  1610 => x"70810651",
  1611 => x"5271802e",
  1612 => x"b13880c6",
  1613 => x"c008ff11",
  1614 => x"545280c6",
  1615 => x"c4087325",
  1616 => x"89387280",
  1617 => x"c6c40cb2",
  1618 => x"e2047110",
  1619 => x"12708429",
  1620 => x"16515288",
  1621 => x"1208802e",
  1622 => x"8938fc51",
  1623 => x"88120852",
  1624 => x"712d80c6",
  1625 => x"c4087053",
  1626 => x"5473802e",
  1627 => x"8a388c15",
  1628 => x"ff155555",
  1629 => x"b2e90482",
  1630 => x"0bbca00c",
  1631 => x"718f06bc",
  1632 => x"9c0c81eb",
  1633 => x"51a9fb2d",
  1634 => x"bc8c0881",
  1635 => x"2a708106",
  1636 => x"51527180",
  1637 => x"2ea73874",
  1638 => x"08852e09",
  1639 => x"81069e38",
  1640 => x"881533ff",
  1641 => x"05527188",
  1642 => x"16347198",
  1643 => x"2b527180",
  1644 => x"25863880",
  1645 => x"0b881634",
  1646 => x"7451aaf2",
  1647 => x"2d81f451",
  1648 => x"a9fb2dbc",
  1649 => x"8c08812a",
  1650 => x"70810651",
  1651 => x"5271802e",
  1652 => x"ab387408",
  1653 => x"852e0981",
  1654 => x"06a23888",
  1655 => x"15338105",
  1656 => x"52718816",
  1657 => x"347181ff",
  1658 => x"068b1633",
  1659 => x"54527272",
  1660 => x"27853872",
  1661 => x"88163474",
  1662 => x"51aaf22d",
  1663 => x"80da51a9",
  1664 => x"fb2dbc8c",
  1665 => x"08812a70",
  1666 => x"81065152",
  1667 => x"71802e81",
  1668 => x"a63880c6",
  1669 => x"bc0880c6",
  1670 => x"c4085553",
  1671 => x"73802e8a",
  1672 => x"388c13ff",
  1673 => x"155553b4",
  1674 => x"9c047208",
  1675 => x"5271822e",
  1676 => x"a6387182",
  1677 => x"26893871",
  1678 => x"812eaa38",
  1679 => x"b5b70471",
  1680 => x"832eb438",
  1681 => x"71842e09",
  1682 => x"810680eb",
  1683 => x"38881308",
  1684 => x"51acbd2d",
  1685 => x"b5b70480",
  1686 => x"c6c40851",
  1687 => x"88130852",
  1688 => x"712db5b7",
  1689 => x"04810b88",
  1690 => x"14082b80",
  1691 => x"c6b00832",
  1692 => x"80c6b00c",
  1693 => x"b58c0488",
  1694 => x"13338105",
  1695 => x"8b143353",
  1696 => x"54717424",
  1697 => x"83388054",
  1698 => x"73881434",
  1699 => x"ab9e2db5",
  1700 => x"b7047508",
  1701 => x"802ea338",
  1702 => x"750851a9",
  1703 => x"fb2dbc8c",
  1704 => x"08810652",
  1705 => x"71802e8c",
  1706 => x"3880c6c4",
  1707 => x"08518416",
  1708 => x"0852712d",
  1709 => x"88165675",
  1710 => x"d9388054",
  1711 => x"800bbca0",
  1712 => x"0c738f06",
  1713 => x"bc9c0ca0",
  1714 => x"527380c6",
  1715 => x"c4082e09",
  1716 => x"81069938",
  1717 => x"80c6c008",
  1718 => x"ff057432",
  1719 => x"70098105",
  1720 => x"7072079f",
  1721 => x"2a917131",
  1722 => x"51515353",
  1723 => x"715182f2",
  1724 => x"2d811454",
  1725 => x"8e7425c4",
  1726 => x"38bc8808",
  1727 => x"5271bc8c",
  1728 => x"0c029805",
  1729 => x"0d040000",
  1730 => x"52657365",
  1731 => x"74000000",
  1732 => x"53617665",
  1733 => x"20736574",
  1734 => x"74696e67",
  1735 => x"73000000",
  1736 => x"5363616e",
  1737 => x"6c696e65",
  1738 => x"73000000",
  1739 => x"4c6f6164",
  1740 => x"20524f4d",
  1741 => x"20100000",
  1742 => x"45786974",
  1743 => x"00000000",
  1744 => x"50432045",
  1745 => x"6e67696e",
  1746 => x"65206d6f",
  1747 => x"64650000",
  1748 => x"54757262",
  1749 => x"6f677261",
  1750 => x"66782031",
  1751 => x"36206d6f",
  1752 => x"64650000",
  1753 => x"56474120",
  1754 => x"2d203331",
  1755 => x"4b487a2c",
  1756 => x"20363048",
  1757 => x"7a000000",
  1758 => x"5456202d",
  1759 => x"20343830",
  1760 => x"692c2036",
  1761 => x"30487a00",
  1762 => x"4261636b",
  1763 => x"00000000",
  1764 => x"46504741",
  1765 => x"50434520",
  1766 => x"43464700",
  1767 => x"496e6974",
  1768 => x"69616c69",
  1769 => x"7a696e67",
  1770 => x"20534420",
  1771 => x"63617264",
  1772 => x"0a000000",
  1773 => x"424f4f54",
  1774 => x"20202020",
  1775 => x"50434500",
  1776 => x"43617264",
  1777 => x"20696e69",
  1778 => x"74206661",
  1779 => x"696c6564",
  1780 => x"0a000000",
  1781 => x"4d425220",
  1782 => x"6661696c",
  1783 => x"0a000000",
  1784 => x"46415431",
  1785 => x"36202020",
  1786 => x"00000000",
  1787 => x"46415433",
  1788 => x"32202020",
  1789 => x"00000000",
  1790 => x"4e6f2070",
  1791 => x"61727469",
  1792 => x"74696f6e",
  1793 => x"20736967",
  1794 => x"0a000000",
  1795 => x"42616420",
  1796 => x"70617274",
  1797 => x"0a000000",
  1798 => x"53444843",
  1799 => x"20657272",
  1800 => x"6f72210a",
  1801 => x"00000000",
  1802 => x"53442069",
  1803 => x"6e69742e",
  1804 => x"2e2e0a00",
  1805 => x"53442063",
  1806 => x"61726420",
  1807 => x"72657365",
  1808 => x"74206661",
  1809 => x"696c6564",
  1810 => x"210a0000",
  1811 => x"57726974",
  1812 => x"65206661",
  1813 => x"696c6564",
  1814 => x"0a000000",
  1815 => x"52656164",
  1816 => x"20666169",
  1817 => x"6c65640a",
  1818 => x"00000000",
  1819 => x"16200000",
  1820 => x"14200000",
  1821 => x"15200000",
  1822 => x"00000002",
  1823 => x"00000002",
  1824 => x"00001b08",
  1825 => x"000004ba",
  1826 => x"00000002",
  1827 => x"00001b10",
  1828 => x"00000379",
  1829 => x"00000003",
  1830 => x"00001ce4",
  1831 => x"00000002",
  1832 => x"00000001",
  1833 => x"00001b20",
  1834 => x"00000001",
  1835 => x"00000003",
  1836 => x"00001cdc",
  1837 => x"00000002",
  1838 => x"00000002",
  1839 => x"00001b2c",
  1840 => x"0000076d",
  1841 => x"00000002",
  1842 => x"00001b38",
  1843 => x"0000155f",
  1844 => x"00000000",
  1845 => x"00000000",
  1846 => x"00000000",
  1847 => x"00001b40",
  1848 => x"00001b50",
  1849 => x"00001b64",
  1850 => x"00001b78",
  1851 => x"0000004d",
  1852 => x"00000741",
  1853 => x"0000002c",
  1854 => x"00000757",
  1855 => x"00000000",
  1856 => x"00000000",
  1857 => x"00000002",
  1858 => x"00001e3c",
  1859 => x"00000542",
  1860 => x"00000002",
  1861 => x"00001e5a",
  1862 => x"00000542",
  1863 => x"00000002",
  1864 => x"00001e78",
  1865 => x"00000542",
  1866 => x"00000002",
  1867 => x"00001e96",
  1868 => x"00000542",
  1869 => x"00000002",
  1870 => x"00001eb4",
  1871 => x"00000542",
  1872 => x"00000002",
  1873 => x"00001ed2",
  1874 => x"00000542",
  1875 => x"00000002",
  1876 => x"00001ef0",
  1877 => x"00000542",
  1878 => x"00000002",
  1879 => x"00001f0e",
  1880 => x"00000542",
  1881 => x"00000002",
  1882 => x"00001f2c",
  1883 => x"00000542",
  1884 => x"00000002",
  1885 => x"00001f4a",
  1886 => x"00000542",
  1887 => x"00000002",
  1888 => x"00001f68",
  1889 => x"00000542",
  1890 => x"00000002",
  1891 => x"00001f86",
  1892 => x"00000542",
  1893 => x"00000002",
  1894 => x"00001fa4",
  1895 => x"00000542",
  1896 => x"00000004",
  1897 => x"00001b88",
  1898 => x"00001c7c",
  1899 => x"00000000",
  1900 => x"00000000",
  1901 => x"000006d5",
  1902 => x"00000000",
  1903 => x"00000000",
  1904 => x"00000000",
  1905 => x"00000000",
  1906 => x"00000000",
  1907 => x"00000000",
  1908 => x"00000000",
  1909 => x"00000000",
  1910 => x"00000000",
  1911 => x"00000000",
  1912 => x"00000000",
  1913 => x"00000000",
  1914 => x"00000000",
  1915 => x"00000000",
  1916 => x"00000000",
  1917 => x"00000000",
  1918 => x"00000000",
  1919 => x"00000000",
  1920 => x"00000000",
  1921 => x"00000000",
  1922 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

