-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bad",
     9 => x"b0080b0b",
    10 => x"0badb408",
    11 => x"0b0b0bad",
    12 => x"b8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"adb80c0b",
    16 => x"0b0badb4",
    17 => x"0c0b0b0b",
    18 => x"adb00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba8c0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"adb070b2",
    57 => x"cc278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8ab30402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"adc00c9f",
    65 => x"0badc40c",
    66 => x"a0717081",
    67 => x"055334ad",
    68 => x"c408ff05",
    69 => x"adc40cad",
    70 => x"c4088025",
    71 => x"eb38adc0",
    72 => x"08ff05ad",
    73 => x"c00cadc0",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0badc0",
    94 => x"08258f38",
    95 => x"82b22dad",
    96 => x"c008ff05",
    97 => x"adc00c82",
    98 => x"f404adc0",
    99 => x"08adc408",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38adc008",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134ad",
   108 => x"c4088105",
   109 => x"adc40cad",
   110 => x"c408519f",
   111 => x"7125e238",
   112 => x"800badc4",
   113 => x"0cadc008",
   114 => x"8105adc0",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"adc40881",
   120 => x"05adc40c",
   121 => x"adc408a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"adc40cad",
   125 => x"c0088105",
   126 => x"adc00c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bad",
   155 => x"c80cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820badc8",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"adc80884",
   167 => x"07adc80c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0bab",
   172 => x"fc0c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cadc808",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f8050d",
   198 => x"b2bc0882",
   199 => x"06aca00b",
   200 => x"80f52d52",
   201 => x"5270802e",
   202 => x"85387181",
   203 => x"0752acac",
   204 => x"0b80f52d",
   205 => x"5170802e",
   206 => x"85387184",
   207 => x"075271ad",
   208 => x"b00c0288",
   209 => x"050d0402",
   210 => x"f4050d74",
   211 => x"708206b2",
   212 => x"bc0cac98",
   213 => x"71810654",
   214 => x"54517188",
   215 => x"1481b72d",
   216 => x"70840651",
   217 => x"70941481",
   218 => x"b72d70ad",
   219 => x"b00c028c",
   220 => x"050d0402",
   221 => x"d4050d7c",
   222 => x"a9c45255",
   223 => x"85f32d99",
   224 => x"db2dadb0",
   225 => x"08802e82",
   226 => x"d0388694",
   227 => x"2dadb008",
   228 => x"538cab2d",
   229 => x"adb00854",
   230 => x"adb00880",
   231 => x"2e82bc38",
   232 => x"840bfec4",
   233 => x"0ca9dc52",
   234 => x"add05192",
   235 => x"bd2dadb0",
   236 => x"08802e80",
   237 => x"ca387482",
   238 => x"2e098106",
   239 => x"a63872ad",
   240 => x"dc0cade0",
   241 => x"5480fd53",
   242 => x"80747084",
   243 => x"05560cff",
   244 => x"13537280",
   245 => x"25f238ad",
   246 => x"dc52add0",
   247 => x"5195a82d",
   248 => x"87ff0474",
   249 => x"812e0981",
   250 => x"069538ad",
   251 => x"dc52add0",
   252 => x"5195822d",
   253 => x"addc0870",
   254 => x"fec00c51",
   255 => x"86c72da9",
   256 => x"e85185f3",
   257 => x"2daa8052",
   258 => x"add05192",
   259 => x"bd2dadb0",
   260 => x"089838aa",
   261 => x"8c5185f3",
   262 => x"2daaa452",
   263 => x"add05192",
   264 => x"bd2dadb0",
   265 => x"08802e81",
   266 => x"b038aab0",
   267 => x"5185f32d",
   268 => x"add40857",
   269 => x"8077595a",
   270 => x"767a2e8b",
   271 => x"38811a78",
   272 => x"812a595a",
   273 => x"77f738f7",
   274 => x"1a5a8077",
   275 => x"25818038",
   276 => x"79527751",
   277 => x"84802dad",
   278 => x"dc52add0",
   279 => x"5195822d",
   280 => x"adb00853",
   281 => x"adb00880",
   282 => x"2e80c938",
   283 => x"addc5b80",
   284 => x"5989a104",
   285 => x"7a708405",
   286 => x"5c087081",
   287 => x"ff067188",
   288 => x"2c7081ff",
   289 => x"0673902c",
   290 => x"7081ff06",
   291 => x"75982afe",
   292 => x"c80cfec8",
   293 => x"0c58fec8",
   294 => x"0c57fec8",
   295 => x"0c841a5a",
   296 => x"53765384",
   297 => x"80772584",
   298 => x"38848053",
   299 => x"727924c4",
   300 => x"3889bf04",
   301 => x"aac05185",
   302 => x"f32d7254",
   303 => x"89db04ad",
   304 => x"d05194d5",
   305 => x"2dfc8017",
   306 => x"81195957",
   307 => x"88ca0482",
   308 => x"0bfec40c",
   309 => x"815489db",
   310 => x"04805473",
   311 => x"adb00c02",
   312 => x"ac050d04",
   313 => x"02f8050d",
   314 => x"a1fe2d81",
   315 => x"f72d8151",
   316 => x"84e52dfe",
   317 => x"c4528172",
   318 => x"0c9fc42d",
   319 => x"9fc42d84",
   320 => x"720c7351",
   321 => x"86f32dac",
   322 => x"8051a3dc",
   323 => x"2d805184",
   324 => x"e52d0288",
   325 => x"050d0402",
   326 => x"fc050d82",
   327 => x"5189e42d",
   328 => x"0284050d",
   329 => x"0402fc05",
   330 => x"0d805189",
   331 => x"e42d0284",
   332 => x"050d0402",
   333 => x"f4050d84",
   334 => x"b85186c7",
   335 => x"2d810bfe",
   336 => x"c40c84b8",
   337 => x"0bfec00c",
   338 => x"840bfec4",
   339 => x"0c830bfe",
   340 => x"cc0c9fdf",
   341 => x"2da1f22d",
   342 => x"9fc42d9f",
   343 => x"c42d81f7",
   344 => x"2d815184",
   345 => x"e52d9fc4",
   346 => x"2d9fc42d",
   347 => x"815184e5",
   348 => x"2d815186",
   349 => x"f32dadb0",
   350 => x"08802e80",
   351 => x"db388051",
   352 => x"84e52dac",
   353 => x"8051a3dc",
   354 => x"2d9ff72d",
   355 => x"a3ec2dad",
   356 => x"b0085386",
   357 => x"942dadb0",
   358 => x"08fec00c",
   359 => x"86942dad",
   360 => x"b008adcc",
   361 => x"082e9c38",
   362 => x"adb008ad",
   363 => x"cc0c8452",
   364 => x"725184e5",
   365 => x"2d9fc42d",
   366 => x"9fc42dff",
   367 => x"12527180",
   368 => x"25ee3872",
   369 => x"802e8938",
   370 => x"8a0bfec4",
   371 => x"0c8b8904",
   372 => x"820bfec4",
   373 => x"0c8b8904",
   374 => x"aad05185",
   375 => x"f32d820b",
   376 => x"fec40c80",
   377 => x"0badb00c",
   378 => x"028c050d",
   379 => x"0402e805",
   380 => x"0d77797b",
   381 => x"58555580",
   382 => x"53727625",
   383 => x"a3387470",
   384 => x"81055680",
   385 => x"f52d7470",
   386 => x"81055680",
   387 => x"f52d5252",
   388 => x"71712e86",
   389 => x"3881518c",
   390 => x"a2048113",
   391 => x"538bf904",
   392 => x"805170ad",
   393 => x"b00c0298",
   394 => x"050d0402",
   395 => x"d8050d80",
   396 => x"0bb1e40c",
   397 => x"addc5280",
   398 => x"519cc32d",
   399 => x"adb00854",
   400 => x"adb0088c",
   401 => x"38aae851",
   402 => x"85f32d73",
   403 => x"5591c604",
   404 => x"8056810b",
   405 => x"b2880c88",
   406 => x"53aaf452",
   407 => x"ae92518b",
   408 => x"ed2dadb0",
   409 => x"08762e09",
   410 => x"81068738",
   411 => x"adb008b2",
   412 => x"880c8853",
   413 => x"ab8052ae",
   414 => x"ae518bed",
   415 => x"2dadb008",
   416 => x"8738adb0",
   417 => x"08b2880c",
   418 => x"b2880880",
   419 => x"2e80f638",
   420 => x"b1a20b80",
   421 => x"f52db1a3",
   422 => x"0b80f52d",
   423 => x"71982b71",
   424 => x"902b07b1",
   425 => x"a40b80f5",
   426 => x"2d70882b",
   427 => x"7207b1a5",
   428 => x"0b80f52d",
   429 => x"7107b1da",
   430 => x"0b80f52d",
   431 => x"b1db0b80",
   432 => x"f52d7188",
   433 => x"2b07535f",
   434 => x"54525a56",
   435 => x"57557381",
   436 => x"abaa2e09",
   437 => x"81068d38",
   438 => x"75519dde",
   439 => x"2dadb008",
   440 => x"568df104",
   441 => x"7382d4d5",
   442 => x"2e8738ab",
   443 => x"8c518eb2",
   444 => x"04addc52",
   445 => x"75519cc3",
   446 => x"2dadb008",
   447 => x"55adb008",
   448 => x"802e83c2",
   449 => x"388853ab",
   450 => x"8052aeae",
   451 => x"518bed2d",
   452 => x"adb00889",
   453 => x"38810bb1",
   454 => x"e40c8eb8",
   455 => x"048853aa",
   456 => x"f452ae92",
   457 => x"518bed2d",
   458 => x"adb00880",
   459 => x"2e8a38ab",
   460 => x"a05185f3",
   461 => x"2d8f9204",
   462 => x"b1da0b80",
   463 => x"f52d5473",
   464 => x"80d52e09",
   465 => x"810680ca",
   466 => x"38b1db0b",
   467 => x"80f52d54",
   468 => x"7381aa2e",
   469 => x"098106ba",
   470 => x"38800bad",
   471 => x"dc0b80f5",
   472 => x"2d565474",
   473 => x"81e92e83",
   474 => x"38815474",
   475 => x"81eb2e8c",
   476 => x"38805573",
   477 => x"752e0981",
   478 => x"0682cb38",
   479 => x"ade70b80",
   480 => x"f52d5574",
   481 => x"8d38ade8",
   482 => x"0b80f52d",
   483 => x"5473822e",
   484 => x"86388055",
   485 => x"91c604ad",
   486 => x"e90b80f5",
   487 => x"2d70b1dc",
   488 => x"0cff05b1",
   489 => x"e00cadea",
   490 => x"0b80f52d",
   491 => x"adeb0b80",
   492 => x"f52d5876",
   493 => x"05778280",
   494 => x"290570b1",
   495 => x"e80cadec",
   496 => x"0b80f52d",
   497 => x"70b1fc0c",
   498 => x"b1e40859",
   499 => x"57587680",
   500 => x"2e81a338",
   501 => x"8853ab80",
   502 => x"52aeae51",
   503 => x"8bed2dad",
   504 => x"b00881e2",
   505 => x"38b1dc08",
   506 => x"70842bb2",
   507 => x"800c70b1",
   508 => x"f80cae81",
   509 => x"0b80f52d",
   510 => x"ae800b80",
   511 => x"f52d7182",
   512 => x"802905ae",
   513 => x"820b80f5",
   514 => x"2d708480",
   515 => x"802912ae",
   516 => x"830b80f5",
   517 => x"2d708180",
   518 => x"0a291270",
   519 => x"b2840cb1",
   520 => x"fc087129",
   521 => x"b1e80805",
   522 => x"70b1ec0c",
   523 => x"ae890b80",
   524 => x"f52dae88",
   525 => x"0b80f52d",
   526 => x"71828029",
   527 => x"05ae8a0b",
   528 => x"80f52d70",
   529 => x"84808029",
   530 => x"12ae8b0b",
   531 => x"80f52d70",
   532 => x"982b81f0",
   533 => x"0a067205",
   534 => x"70b1f00c",
   535 => x"fe117e29",
   536 => x"7705b1f4",
   537 => x"0c525952",
   538 => x"43545e51",
   539 => x"5259525d",
   540 => x"57595791",
   541 => x"c404adee",
   542 => x"0b80f52d",
   543 => x"aded0b80",
   544 => x"f52d7182",
   545 => x"80290570",
   546 => x"b2800c70",
   547 => x"a02983ff",
   548 => x"0570892a",
   549 => x"70b1f80c",
   550 => x"adf30b80",
   551 => x"f52dadf2",
   552 => x"0b80f52d",
   553 => x"71828029",
   554 => x"0570b284",
   555 => x"0c7b7129",
   556 => x"1e70b1f4",
   557 => x"0c7db1f0",
   558 => x"0c7305b1",
   559 => x"ec0c555e",
   560 => x"51515555",
   561 => x"815574ad",
   562 => x"b00c02a8",
   563 => x"050d0402",
   564 => x"ec050d76",
   565 => x"70872c71",
   566 => x"80ff0655",
   567 => x"5654b1e4",
   568 => x"088a3873",
   569 => x"882c7481",
   570 => x"ff065455",
   571 => x"addc52b1",
   572 => x"e8081551",
   573 => x"9cc32dad",
   574 => x"b00854ad",
   575 => x"b008802e",
   576 => x"b338b1e4",
   577 => x"08802e98",
   578 => x"38728429",
   579 => x"addc0570",
   580 => x"0852539d",
   581 => x"de2dadb0",
   582 => x"08f00a06",
   583 => x"5392b204",
   584 => x"7210addc",
   585 => x"057080e0",
   586 => x"2d52539e",
   587 => x"8e2dadb0",
   588 => x"08537254",
   589 => x"73adb00c",
   590 => x"0294050d",
   591 => x"0402c805",
   592 => x"0d7f615f",
   593 => x"5b800bb1",
   594 => x"f008b1f4",
   595 => x"08595d56",
   596 => x"b1e40876",
   597 => x"2e8a38b1",
   598 => x"dc08842b",
   599 => x"5892e604",
   600 => x"b1f80884",
   601 => x"2b588059",
   602 => x"78782781",
   603 => x"a938788f",
   604 => x"06a01757",
   605 => x"54738f38",
   606 => x"addc5276",
   607 => x"51811757",
   608 => x"9cc32dad",
   609 => x"dc568076",
   610 => x"80f52d56",
   611 => x"5474742e",
   612 => x"83388154",
   613 => x"7481e52e",
   614 => x"80f63881",
   615 => x"70750655",
   616 => x"5d73802e",
   617 => x"80ea388b",
   618 => x"1680f52d",
   619 => x"98065a79",
   620 => x"80de388b",
   621 => x"537d5275",
   622 => x"518bed2d",
   623 => x"adb00880",
   624 => x"cf389c16",
   625 => x"08519dde",
   626 => x"2dadb008",
   627 => x"841c0c9a",
   628 => x"1680e02d",
   629 => x"519e8e2d",
   630 => x"adb008ad",
   631 => x"b008881d",
   632 => x"0cadb008",
   633 => x"5555b1e4",
   634 => x"08802e98",
   635 => x"38941680",
   636 => x"e02d519e",
   637 => x"8e2dadb0",
   638 => x"08902b83",
   639 => x"fff00a06",
   640 => x"70165154",
   641 => x"73881c0c",
   642 => x"797b0c7c",
   643 => x"5494cc04",
   644 => x"81195992",
   645 => x"e804b1e4",
   646 => x"08802eae",
   647 => x"387b5191",
   648 => x"cf2dadb0",
   649 => x"08adb008",
   650 => x"80ffffff",
   651 => x"f806555c",
   652 => x"7380ffff",
   653 => x"fff82e92",
   654 => x"38adb008",
   655 => x"fe05b1dc",
   656 => x"0829b1ec",
   657 => x"08055792",
   658 => x"e6048054",
   659 => x"73adb00c",
   660 => x"02b8050d",
   661 => x"0402f405",
   662 => x"0d747008",
   663 => x"8105710c",
   664 => x"7008b1e0",
   665 => x"08065353",
   666 => x"718e3888",
   667 => x"13085191",
   668 => x"cf2dadb0",
   669 => x"0888140c",
   670 => x"810badb0",
   671 => x"0c028c05",
   672 => x"0d0402f0",
   673 => x"050d7588",
   674 => x"1108fe05",
   675 => x"b1dc0829",
   676 => x"b1ec0811",
   677 => x"7208b1e0",
   678 => x"08060579",
   679 => x"55535454",
   680 => x"9cc32d02",
   681 => x"90050d04",
   682 => x"02f0050d",
   683 => x"75881108",
   684 => x"fe05b1dc",
   685 => x"0829b1ec",
   686 => x"08117208",
   687 => x"b1e00806",
   688 => x"05795553",
   689 => x"54549b83",
   690 => x"2d029005",
   691 => x"0d0402f4",
   692 => x"050dd452",
   693 => x"81ff720c",
   694 => x"71085381",
   695 => x"ff720c72",
   696 => x"882b83fe",
   697 => x"80067208",
   698 => x"7081ff06",
   699 => x"51525381",
   700 => x"ff720c72",
   701 => x"7107882b",
   702 => x"72087081",
   703 => x"ff065152",
   704 => x"5381ff72",
   705 => x"0c727107",
   706 => x"882b7208",
   707 => x"7081ff06",
   708 => x"7207adb0",
   709 => x"0c525302",
   710 => x"8c050d04",
   711 => x"02f4050d",
   712 => x"74767181",
   713 => x"ff06d40c",
   714 => x"5353b28c",
   715 => x"08853871",
   716 => x"892b5271",
   717 => x"982ad40c",
   718 => x"71902a70",
   719 => x"81ff06d4",
   720 => x"0c517188",
   721 => x"2a7081ff",
   722 => x"06d40c51",
   723 => x"7181ff06",
   724 => x"d40c7290",
   725 => x"2a7081ff",
   726 => x"06d40c51",
   727 => x"d4087081",
   728 => x"ff065151",
   729 => x"82b8bf52",
   730 => x"7081ff2e",
   731 => x"09810694",
   732 => x"3881ff0b",
   733 => x"d40cd408",
   734 => x"7081ff06",
   735 => x"ff145451",
   736 => x"5171e538",
   737 => x"70adb00c",
   738 => x"028c050d",
   739 => x"0402fc05",
   740 => x"0d81c751",
   741 => x"81ff0bd4",
   742 => x"0cff1151",
   743 => x"708025f4",
   744 => x"38028405",
   745 => x"0d0402f0",
   746 => x"050d978d",
   747 => x"2d8fcf53",
   748 => x"805287fc",
   749 => x"80f75196",
   750 => x"9c2dadb0",
   751 => x"0854adb0",
   752 => x"08812e09",
   753 => x"8106a338",
   754 => x"81ff0bd4",
   755 => x"0c820a52",
   756 => x"849c80e9",
   757 => x"51969c2d",
   758 => x"adb0088b",
   759 => x"3881ff0b",
   760 => x"d40c7353",
   761 => x"97f00497",
   762 => x"8d2dff13",
   763 => x"5372c138",
   764 => x"72adb00c",
   765 => x"0290050d",
   766 => x"0402f405",
   767 => x"0d81ff0b",
   768 => x"d40c9353",
   769 => x"805287fc",
   770 => x"80c15196",
   771 => x"9c2dadb0",
   772 => x"088b3881",
   773 => x"ff0bd40c",
   774 => x"815398a6",
   775 => x"04978d2d",
   776 => x"ff135372",
   777 => x"df3872ad",
   778 => x"b00c028c",
   779 => x"050d0402",
   780 => x"f0050d97",
   781 => x"8d2d83aa",
   782 => x"52849c80",
   783 => x"c851969c",
   784 => x"2dadb008",
   785 => x"812e0981",
   786 => x"06923895",
   787 => x"ce2dadb0",
   788 => x"0883ffff",
   789 => x"06537283",
   790 => x"aa2e9738",
   791 => x"97f92d98",
   792 => x"ed048154",
   793 => x"99d204ab",
   794 => x"ac5185f3",
   795 => x"2d805499",
   796 => x"d20481ff",
   797 => x"0bd40cb1",
   798 => x"5397a62d",
   799 => x"adb00880",
   800 => x"2e80c038",
   801 => x"805287fc",
   802 => x"80fa5196",
   803 => x"9c2dadb0",
   804 => x"08b13881",
   805 => x"ff0bd40c",
   806 => x"d4085381",
   807 => x"ff0bd40c",
   808 => x"81ff0bd4",
   809 => x"0c81ff0b",
   810 => x"d40c81ff",
   811 => x"0bd40c72",
   812 => x"862a7081",
   813 => x"06adb008",
   814 => x"56515372",
   815 => x"802e9338",
   816 => x"98e20472",
   817 => x"822eff9f",
   818 => x"38ff1353",
   819 => x"72ffaa38",
   820 => x"725473ad",
   821 => x"b00c0290",
   822 => x"050d0402",
   823 => x"f0050d81",
   824 => x"0bb28c0c",
   825 => x"8454d008",
   826 => x"708f2a70",
   827 => x"81065151",
   828 => x"5372f338",
   829 => x"72d00c97",
   830 => x"8d2dabbc",
   831 => x"5185f32d",
   832 => x"d008708f",
   833 => x"2a708106",
   834 => x"51515372",
   835 => x"f338810b",
   836 => x"d00cb153",
   837 => x"805284d4",
   838 => x"80c05196",
   839 => x"9c2dadb0",
   840 => x"08812ea1",
   841 => x"3872822e",
   842 => x"0981068c",
   843 => x"38abc851",
   844 => x"85f32d80",
   845 => x"539afa04",
   846 => x"ff135372",
   847 => x"d738ff14",
   848 => x"5473ffa2",
   849 => x"3898af2d",
   850 => x"adb008b2",
   851 => x"8c0cadb0",
   852 => x"088b3881",
   853 => x"5287fc80",
   854 => x"d051969c",
   855 => x"2d81ff0b",
   856 => x"d40cd008",
   857 => x"708f2a70",
   858 => x"81065151",
   859 => x"5372f338",
   860 => x"72d00c81",
   861 => x"ff0bd40c",
   862 => x"815372ad",
   863 => x"b00c0290",
   864 => x"050d0402",
   865 => x"e8050d78",
   866 => x"5681ff0b",
   867 => x"d40cd008",
   868 => x"708f2a70",
   869 => x"81065151",
   870 => x"5372f338",
   871 => x"82810bd0",
   872 => x"0c81ff0b",
   873 => x"d40c7752",
   874 => x"87fc80d8",
   875 => x"51969c2d",
   876 => x"adb00880",
   877 => x"2e8c38ab",
   878 => x"e05185f3",
   879 => x"2d81539c",
   880 => x"ba0481ff",
   881 => x"0bd40c81",
   882 => x"fe0bd40c",
   883 => x"80ff5575",
   884 => x"70840557",
   885 => x"0870982a",
   886 => x"d40c7090",
   887 => x"2c7081ff",
   888 => x"06d40c54",
   889 => x"70882c70",
   890 => x"81ff06d4",
   891 => x"0c547081",
   892 => x"ff06d40c",
   893 => x"54ff1555",
   894 => x"748025d3",
   895 => x"3881ff0b",
   896 => x"d40c81ff",
   897 => x"0bd40c81",
   898 => x"ff0bd40c",
   899 => x"868da054",
   900 => x"81ff0bd4",
   901 => x"0cd40881",
   902 => x"ff065574",
   903 => x"8738ff14",
   904 => x"5473ed38",
   905 => x"81ff0bd4",
   906 => x"0cd00870",
   907 => x"8f2a7081",
   908 => x"06515153",
   909 => x"72f33872",
   910 => x"d00c72ad",
   911 => x"b00c0298",
   912 => x"050d0402",
   913 => x"e8050d78",
   914 => x"55805681",
   915 => x"ff0bd40c",
   916 => x"d008708f",
   917 => x"2a708106",
   918 => x"51515372",
   919 => x"f3388281",
   920 => x"0bd00c81",
   921 => x"ff0bd40c",
   922 => x"775287fc",
   923 => x"80d15196",
   924 => x"9c2d80db",
   925 => x"c6df54ad",
   926 => x"b008802e",
   927 => x"8a38aac0",
   928 => x"5185f32d",
   929 => x"9dd50481",
   930 => x"ff0bd40c",
   931 => x"d4087081",
   932 => x"ff065153",
   933 => x"7281fe2e",
   934 => x"0981069d",
   935 => x"3880ff53",
   936 => x"95ce2dad",
   937 => x"b0087570",
   938 => x"8405570c",
   939 => x"ff135372",
   940 => x"8025ed38",
   941 => x"81569dbf",
   942 => x"04ff1454",
   943 => x"73c93881",
   944 => x"ff0bd40c",
   945 => x"d008708f",
   946 => x"2a708106",
   947 => x"51515372",
   948 => x"f33872d0",
   949 => x"0c75adb0",
   950 => x"0c029805",
   951 => x"0d0402f4",
   952 => x"050d7470",
   953 => x"882a83fe",
   954 => x"80067072",
   955 => x"982a0772",
   956 => x"882b87fc",
   957 => x"80800673",
   958 => x"982b81f0",
   959 => x"0a067173",
   960 => x"0707adb0",
   961 => x"0c565153",
   962 => x"51028c05",
   963 => x"0d0402f8",
   964 => x"050d028e",
   965 => x"0580f52d",
   966 => x"74882b07",
   967 => x"7083ffff",
   968 => x"06adb00c",
   969 => x"51028805",
   970 => x"0d0402fc",
   971 => x"050d7251",
   972 => x"80710c80",
   973 => x"0b84120c",
   974 => x"0284050d",
   975 => x"0402f005",
   976 => x"0d757008",
   977 => x"84120853",
   978 => x"5353ff54",
   979 => x"71712ea8",
   980 => x"38a1f82d",
   981 => x"84130870",
   982 => x"84291488",
   983 => x"11700870",
   984 => x"81ff0684",
   985 => x"18088111",
   986 => x"8706841a",
   987 => x"0c535155",
   988 => x"515151a1",
   989 => x"f22d7154",
   990 => x"73adb00c",
   991 => x"0290050d",
   992 => x"0402f805",
   993 => x"0da1f82d",
   994 => x"e008708b",
   995 => x"2a708106",
   996 => x"51525270",
   997 => x"802e9d38",
   998 => x"b2900870",
   999 => x"8429b298",
  1000 => x"057381ff",
  1001 => x"06710c51",
  1002 => x"51b29008",
  1003 => x"81118706",
  1004 => x"b2900c51",
  1005 => x"800bb2b8",
  1006 => x"0ca1eb2d",
  1007 => x"a1f22d02",
  1008 => x"88050d04",
  1009 => x"02fc050d",
  1010 => x"a1f82d81",
  1011 => x"0bb2b80c",
  1012 => x"a1f22db2",
  1013 => x"b8085170",
  1014 => x"fa380284",
  1015 => x"050d0402",
  1016 => x"fc050db2",
  1017 => x"90519eaa",
  1018 => x"2d9f8151",
  1019 => x"a1e72da1",
  1020 => x"912d0284",
  1021 => x"050d0402",
  1022 => x"f4050da0",
  1023 => x"f904adb0",
  1024 => x"0881f02e",
  1025 => x"09810689",
  1026 => x"38810bad",
  1027 => x"a40ca0f9",
  1028 => x"04adb008",
  1029 => x"81e02e09",
  1030 => x"81068938",
  1031 => x"810bada8",
  1032 => x"0ca0f904",
  1033 => x"adb00852",
  1034 => x"ada80880",
  1035 => x"2e8838ad",
  1036 => x"b0088180",
  1037 => x"05527184",
  1038 => x"2c728f06",
  1039 => x"5353ada4",
  1040 => x"08802e99",
  1041 => x"38728429",
  1042 => x"ace40572",
  1043 => x"1381712b",
  1044 => x"70097308",
  1045 => x"06730c51",
  1046 => x"5353a0ef",
  1047 => x"04728429",
  1048 => x"ace40572",
  1049 => x"1383712b",
  1050 => x"72080772",
  1051 => x"0c535380",
  1052 => x"0bada80c",
  1053 => x"800bada4",
  1054 => x"0cb29051",
  1055 => x"9ebd2dad",
  1056 => x"b008ff24",
  1057 => x"fef83880",
  1058 => x"0badb00c",
  1059 => x"028c050d",
  1060 => x"0402f805",
  1061 => x"0dace452",
  1062 => x"8f518072",
  1063 => x"70840554",
  1064 => x"0cff1151",
  1065 => x"708025f2",
  1066 => x"38028805",
  1067 => x"0d0402f0",
  1068 => x"050d7551",
  1069 => x"a1f82d70",
  1070 => x"822cfc06",
  1071 => x"ace41172",
  1072 => x"109e0671",
  1073 => x"0870722a",
  1074 => x"70830682",
  1075 => x"742b7009",
  1076 => x"7406760c",
  1077 => x"54515657",
  1078 => x"535153a1",
  1079 => x"f22d71ad",
  1080 => x"b00c0290",
  1081 => x"050d0471",
  1082 => x"980c04ff",
  1083 => x"b008adb0",
  1084 => x"0c04810b",
  1085 => x"ffb00c04",
  1086 => x"800bffb0",
  1087 => x"0c0402fc",
  1088 => x"050d800b",
  1089 => x"adac0c80",
  1090 => x"5184e52d",
  1091 => x"0284050d",
  1092 => x"0402ec05",
  1093 => x"0d765480",
  1094 => x"52870b88",
  1095 => x"1580f52d",
  1096 => x"56537472",
  1097 => x"248338a0",
  1098 => x"53725182",
  1099 => x"ee2d8112",
  1100 => x"8b1580f5",
  1101 => x"2d545272",
  1102 => x"7225de38",
  1103 => x"0294050d",
  1104 => x"0402f005",
  1105 => x"0db2c008",
  1106 => x"5481f72d",
  1107 => x"800bb2c4",
  1108 => x"0c730880",
  1109 => x"2e818038",
  1110 => x"820badc4",
  1111 => x"0cb2c408",
  1112 => x"8f06adc0",
  1113 => x"0c730852",
  1114 => x"71832e96",
  1115 => x"38718326",
  1116 => x"89387181",
  1117 => x"2eaf38a3",
  1118 => x"c2047185",
  1119 => x"2e9f38a3",
  1120 => x"c2048814",
  1121 => x"80f52d84",
  1122 => x"1508abf0",
  1123 => x"53545285",
  1124 => x"f32d7184",
  1125 => x"29137008",
  1126 => x"5252a3c6",
  1127 => x"047351a2",
  1128 => x"912da3c2",
  1129 => x"04b2bc08",
  1130 => x"8815082c",
  1131 => x"70810651",
  1132 => x"5271802e",
  1133 => x"8738abf4",
  1134 => x"51a3bf04",
  1135 => x"abf85185",
  1136 => x"f32d8414",
  1137 => x"085185f3",
  1138 => x"2db2c408",
  1139 => x"8105b2c4",
  1140 => x"0c8c1454",
  1141 => x"a2d10402",
  1142 => x"90050d04",
  1143 => x"71b2c00c",
  1144 => x"a2c12db2",
  1145 => x"c408ff05",
  1146 => x"b2c80c04",
  1147 => x"02ec050d",
  1148 => x"b2c00855",
  1149 => x"80f851a1",
  1150 => x"ae2dadb0",
  1151 => x"08812a70",
  1152 => x"81065152",
  1153 => x"719b3887",
  1154 => x"51a1ae2d",
  1155 => x"adb00881",
  1156 => x"2a708106",
  1157 => x"51527180",
  1158 => x"2eb138a4",
  1159 => x"a1049ff7",
  1160 => x"2d8751a1",
  1161 => x"ae2dadb0",
  1162 => x"08f438a4",
  1163 => x"b1049ff7",
  1164 => x"2d80f851",
  1165 => x"a1ae2dad",
  1166 => x"b008f338",
  1167 => x"adac0881",
  1168 => x"3270adac",
  1169 => x"0c705252",
  1170 => x"84e52dad",
  1171 => x"ac08a238",
  1172 => x"80da51a1",
  1173 => x"ae2d81f5",
  1174 => x"51a1ae2d",
  1175 => x"81f251a1",
  1176 => x"ae2d81eb",
  1177 => x"51a1ae2d",
  1178 => x"81f451a1",
  1179 => x"ae2da8b5",
  1180 => x"0481f551",
  1181 => x"a1ae2dad",
  1182 => x"b008812a",
  1183 => x"70810651",
  1184 => x"5271802e",
  1185 => x"8f38b2c8",
  1186 => x"08527180",
  1187 => x"2e8638ff",
  1188 => x"12b2c80c",
  1189 => x"81f251a1",
  1190 => x"ae2dadb0",
  1191 => x"08812a70",
  1192 => x"81065152",
  1193 => x"71802e95",
  1194 => x"38b2c408",
  1195 => x"ff05b2c8",
  1196 => x"08545272",
  1197 => x"72258638",
  1198 => x"8113b2c8",
  1199 => x"0cb2c808",
  1200 => x"70535473",
  1201 => x"802e8a38",
  1202 => x"8c15ff15",
  1203 => x"5555a5c3",
  1204 => x"04820bad",
  1205 => x"c40c718f",
  1206 => x"06adc00c",
  1207 => x"81eb51a1",
  1208 => x"ae2dadb0",
  1209 => x"08812a70",
  1210 => x"81065152",
  1211 => x"71802ead",
  1212 => x"38740885",
  1213 => x"2e098106",
  1214 => x"a4388815",
  1215 => x"80f52dff",
  1216 => x"05527188",
  1217 => x"1681b72d",
  1218 => x"71982b52",
  1219 => x"71802588",
  1220 => x"38800b88",
  1221 => x"1681b72d",
  1222 => x"7451a291",
  1223 => x"2d81f451",
  1224 => x"a1ae2dad",
  1225 => x"b008812a",
  1226 => x"70810651",
  1227 => x"5271802e",
  1228 => x"b3387408",
  1229 => x"852e0981",
  1230 => x"06aa3888",
  1231 => x"1580f52d",
  1232 => x"81055271",
  1233 => x"881681b7",
  1234 => x"2d7181ff",
  1235 => x"068b1680",
  1236 => x"f52d5452",
  1237 => x"72722787",
  1238 => x"38728816",
  1239 => x"81b72d74",
  1240 => x"51a2912d",
  1241 => x"80da51a1",
  1242 => x"ae2dadb0",
  1243 => x"08812a70",
  1244 => x"81065152",
  1245 => x"71802e80",
  1246 => x"fb38b2c0",
  1247 => x"08b2c808",
  1248 => x"55537380",
  1249 => x"2e8a388c",
  1250 => x"13ff1555",
  1251 => x"53a78204",
  1252 => x"72085271",
  1253 => x"822ea638",
  1254 => x"71822689",
  1255 => x"3871812e",
  1256 => x"a538a7f4",
  1257 => x"0471832e",
  1258 => x"ad387184",
  1259 => x"2e098106",
  1260 => x"80c23888",
  1261 => x"130851a3",
  1262 => x"dc2da7f4",
  1263 => x"04881308",
  1264 => x"52712da7",
  1265 => x"f404810b",
  1266 => x"8814082b",
  1267 => x"b2bc0832",
  1268 => x"b2bc0ca7",
  1269 => x"f1048813",
  1270 => x"80f52d81",
  1271 => x"058b1480",
  1272 => x"f52d5354",
  1273 => x"71742483",
  1274 => x"38805473",
  1275 => x"881481b7",
  1276 => x"2da2c12d",
  1277 => x"8054800b",
  1278 => x"adc40c73",
  1279 => x"8f06adc0",
  1280 => x"0ca05273",
  1281 => x"b2c8082e",
  1282 => x"09810698",
  1283 => x"38b2c408",
  1284 => x"ff057432",
  1285 => x"70098105",
  1286 => x"7072079f",
  1287 => x"2a917131",
  1288 => x"51515353",
  1289 => x"715182ee",
  1290 => x"2d811454",
  1291 => x"8e7425c6",
  1292 => x"38adac08",
  1293 => x"5271adb0",
  1294 => x"0c029405",
  1295 => x"0d040000",
  1296 => x"00ffffff",
  1297 => x"ff00ffff",
  1298 => x"ffff00ff",
  1299 => x"ffffff00",
  1300 => x"52657365",
  1301 => x"74000000",
  1302 => x"53617665",
  1303 => x"20616e64",
  1304 => x"20526573",
  1305 => x"65740000",
  1306 => x"5363616e",
  1307 => x"6c696e65",
  1308 => x"73000000",
  1309 => x"45786974",
  1310 => x"00000000",
  1311 => x"50432045",
  1312 => x"6e67696e",
  1313 => x"65206d6f",
  1314 => x"64650000",
  1315 => x"54757262",
  1316 => x"6f677261",
  1317 => x"66782031",
  1318 => x"36206d6f",
  1319 => x"64650000",
  1320 => x"56474120",
  1321 => x"2d203331",
  1322 => x"4b487a2c",
  1323 => x"20363048",
  1324 => x"7a000000",
  1325 => x"5456202d",
  1326 => x"20343830",
  1327 => x"692c2036",
  1328 => x"30487a00",
  1329 => x"496e6974",
  1330 => x"69616c69",
  1331 => x"7a696e67",
  1332 => x"20534420",
  1333 => x"63617264",
  1334 => x"0a000000",
  1335 => x"46504741",
  1336 => x"50434520",
  1337 => x"43464700",
  1338 => x"54727969",
  1339 => x"6e67204d",
  1340 => x"53583342",
  1341 => x"494f532e",
  1342 => x"5359530a",
  1343 => x"00000000",
  1344 => x"4d535833",
  1345 => x"42494f53",
  1346 => x"53595300",
  1347 => x"54727969",
  1348 => x"6e672042",
  1349 => x"494f535f",
  1350 => x"4d32502e",
  1351 => x"524f4d0a",
  1352 => x"00000000",
  1353 => x"42494f53",
  1354 => x"5f4d3250",
  1355 => x"524f4d00",
  1356 => x"4c6f6164",
  1357 => x"696e6720",
  1358 => x"42494f53",
  1359 => x"0a000000",
  1360 => x"52656164",
  1361 => x"20666169",
  1362 => x"6c65640a",
  1363 => x"00000000",
  1364 => x"4c6f6164",
  1365 => x"696e6720",
  1366 => x"42494f53",
  1367 => x"20666169",
  1368 => x"6c65640a",
  1369 => x"00000000",
  1370 => x"4d425220",
  1371 => x"6661696c",
  1372 => x"0a000000",
  1373 => x"46415431",
  1374 => x"36202020",
  1375 => x"00000000",
  1376 => x"46415433",
  1377 => x"32202020",
  1378 => x"00000000",
  1379 => x"4e6f2070",
  1380 => x"61727469",
  1381 => x"74696f6e",
  1382 => x"20736967",
  1383 => x"0a000000",
  1384 => x"42616420",
  1385 => x"70617274",
  1386 => x"0a000000",
  1387 => x"53444843",
  1388 => x"20657272",
  1389 => x"6f72210a",
  1390 => x"00000000",
  1391 => x"53442069",
  1392 => x"6e69742e",
  1393 => x"2e2e0a00",
  1394 => x"53442063",
  1395 => x"61726420",
  1396 => x"72657365",
  1397 => x"74206661",
  1398 => x"696c6564",
  1399 => x"210a0000",
  1400 => x"57726974",
  1401 => x"65206661",
  1402 => x"696c6564",
  1403 => x"0a000000",
  1404 => x"16200000",
  1405 => x"14200000",
  1406 => x"15200000",
  1407 => x"00000002",
  1408 => x"00000002",
  1409 => x"00001450",
  1410 => x"00000525",
  1411 => x"00000002",
  1412 => x"00001458",
  1413 => x"00000517",
  1414 => x"00000003",
  1415 => x"0000165c",
  1416 => x"00000002",
  1417 => x"00000001",
  1418 => x"00001468",
  1419 => x"0000000b",
  1420 => x"00000003",
  1421 => x"00001654",
  1422 => x"00000002",
  1423 => x"00000002",
  1424 => x"00001474",
  1425 => x"000010fe",
  1426 => x"00000000",
  1427 => x"00000000",
  1428 => x"00000000",
  1429 => x"0000147c",
  1430 => x"0000148c",
  1431 => x"000014a0",
  1432 => x"000014b4",
  1433 => x"00000000",
  1434 => x"00000000",
  1435 => x"00000000",
  1436 => x"00000000",
  1437 => x"00000000",
  1438 => x"00000000",
  1439 => x"00000000",
  1440 => x"00000000",
  1441 => x"00000000",
  1442 => x"00000000",
  1443 => x"00000000",
  1444 => x"00000000",
  1445 => x"00000000",
  1446 => x"00000000",
  1447 => x"00000000",
  1448 => x"00000000",
  1449 => x"00000000",
  1450 => x"00000000",
  1451 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

