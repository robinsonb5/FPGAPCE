-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb6",
     9 => x"c8080b0b",
    10 => x"0bb6cc08",
    11 => x"0b0b0bb6",
    12 => x"d0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b6d00c0b",
    16 => x"0b0bb6cc",
    17 => x"0c0b0b0b",
    18 => x"b6c80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb0b0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b6c870bd",
    57 => x"c4278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8d950402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b6d80c9f",
    65 => x"0bb6dc0c",
    66 => x"a0717081",
    67 => x"055334b6",
    68 => x"dc08ff05",
    69 => x"b6dc0cb6",
    70 => x"dc088025",
    71 => x"eb38b6d8",
    72 => x"08ff05b6",
    73 => x"d80cb6d8",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb6d8",
    94 => x"08258f38",
    95 => x"82b22db6",
    96 => x"d808ff05",
    97 => x"b6d80c82",
    98 => x"f404b6d8",
    99 => x"08b6dc08",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b6d808",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b6",
   108 => x"dc088105",
   109 => x"b6dc0cb6",
   110 => x"dc08519f",
   111 => x"7125e238",
   112 => x"800bb6dc",
   113 => x"0cb6d808",
   114 => x"8105b6d8",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b6dc0881",
   120 => x"05b6dc0c",
   121 => x"b6dc08a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b6dc0cb6",
   125 => x"d8088105",
   126 => x"b6d80c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb6",
   155 => x"e00cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb6e0",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b6e00884",
   167 => x"07b6e00c",
   168 => x"5573842b",
   169 => x"87e87125",
   170 => x"83713170",
   171 => x"0b0b0bb3",
   172 => x"b80c8171",
   173 => x"2bf6880c",
   174 => x"fea413ff",
   175 => x"122c7888",
   176 => x"29ff9405",
   177 => x"70812cb6",
   178 => x"e0085258",
   179 => x"52555152",
   180 => x"5476802e",
   181 => x"85387081",
   182 => x"075170f6",
   183 => x"940c7109",
   184 => x"8105f680",
   185 => x"0c720981",
   186 => x"05f6840c",
   187 => x"0294050d",
   188 => x"0402f405",
   189 => x"0d745372",
   190 => x"70810554",
   191 => x"80f52d52",
   192 => x"71802e89",
   193 => x"38715182",
   194 => x"ee2d85f7",
   195 => x"04028c05",
   196 => x"0d0402f4",
   197 => x"050d7470",
   198 => x"8206bda8",
   199 => x"0cb3d471",
   200 => x"81065454",
   201 => x"51718814",
   202 => x"81b72d70",
   203 => x"822a7081",
   204 => x"06515170",
   205 => x"941481b7",
   206 => x"2d70b6c8",
   207 => x"0c028c05",
   208 => x"0d0402f8",
   209 => x"050db1c8",
   210 => x"52b6e451",
   211 => x"96b32db6",
   212 => x"c808802e",
   213 => x"9d38b8c8",
   214 => x"52b6e451",
   215 => x"98e92db8",
   216 => x"c808b6f0",
   217 => x"0cb8c808",
   218 => x"fec00cb8",
   219 => x"c8085186",
   220 => x"922d0288",
   221 => x"050d0402",
   222 => x"f0050db1",
   223 => x"c852b6e4",
   224 => x"5196b32d",
   225 => x"b6c80880",
   226 => x"2ea538b6",
   227 => x"f008b8c8",
   228 => x"0cb8cc54",
   229 => x"80fd5380",
   230 => x"74708405",
   231 => x"560cff13",
   232 => x"53728025",
   233 => x"f238b8c8",
   234 => x"52b6e451",
   235 => x"998f2d02",
   236 => x"90050d04",
   237 => x"02d8050d",
   238 => x"810bfec4",
   239 => x"0c840bfe",
   240 => x"c40c7b52",
   241 => x"b6e45196",
   242 => x"b32db6c8",
   243 => x"0853b6c8",
   244 => x"08802e81",
   245 => x"d538b6e8",
   246 => x"0856800b",
   247 => x"ff175859",
   248 => x"76792e8b",
   249 => x"38811977",
   250 => x"812a5859",
   251 => x"76f738f7",
   252 => x"19769fff",
   253 => x"06545972",
   254 => x"802e8b38",
   255 => x"fc8016b6",
   256 => x"e4525698",
   257 => x"bc2db6f0",
   258 => x"08f70670",
   259 => x"b6f00c53",
   260 => x"75b08080",
   261 => x"2e098106",
   262 => x"87387288",
   263 => x"07b6f00c",
   264 => x"b6f008fe",
   265 => x"c00c8076",
   266 => x"2580fa38",
   267 => x"78527651",
   268 => x"84802db8",
   269 => x"c852b6e4",
   270 => x"5198e92d",
   271 => x"b6c80853",
   272 => x"b6c80880",
   273 => x"2e80c838",
   274 => x"b8c85a80",
   275 => x"5888fc04",
   276 => x"79708405",
   277 => x"5b087083",
   278 => x"fe800671",
   279 => x"882b83fe",
   280 => x"80067188",
   281 => x"2a077288",
   282 => x"2a83fe80",
   283 => x"0673982a",
   284 => x"07fec80c",
   285 => x"fec80c56",
   286 => x"84195953",
   287 => x"75538480",
   288 => x"76258438",
   289 => x"84805372",
   290 => x"7824c538",
   291 => x"899504b1",
   292 => x"d45189ad",
   293 => x"04b6e451",
   294 => x"98bc2dfc",
   295 => x"80168118",
   296 => x"585688a6",
   297 => x"04815389",
   298 => x"b004b1e4",
   299 => x"5185f12d",
   300 => x"72b6c80c",
   301 => x"02a8050d",
   302 => x"0402fc05",
   303 => x"0da5fd2d",
   304 => x"fec45181",
   305 => x"710c8271",
   306 => x"0c028405",
   307 => x"0d0402f4",
   308 => x"050d7410",
   309 => x"15708429",
   310 => x"b4c80570",
   311 => x"08555152",
   312 => x"72802e90",
   313 => x"387280f5",
   314 => x"2d527180",
   315 => x"2e863872",
   316 => x"5187b42d",
   317 => x"b3bc51a7",
   318 => x"db2da5fd",
   319 => x"2d805184",
   320 => x"e52d028c",
   321 => x"050d0402",
   322 => x"e8050d80",
   323 => x"70565675",
   324 => x"b5f80825",
   325 => x"af38bcd4",
   326 => x"08762ea8",
   327 => x"38745195",
   328 => x"de2db6c8",
   329 => x"08098105",
   330 => x"70b6c808",
   331 => x"079f2a77",
   332 => x"05811757",
   333 => x"575275b5",
   334 => x"f8082588",
   335 => x"38bcd408",
   336 => x"7526da38",
   337 => x"805674bc",
   338 => x"d4082780",
   339 => x"d0387451",
   340 => x"95de2d75",
   341 => x"842b52b6",
   342 => x"c808802e",
   343 => x"ae38b6f8",
   344 => x"128117b6",
   345 => x"c8085657",
   346 => x"528a5373",
   347 => x"70810555",
   348 => x"80f52d72",
   349 => x"70810554",
   350 => x"81b72dff",
   351 => x"13537280",
   352 => x"25e93880",
   353 => x"7281b72d",
   354 => x"8b9404b6",
   355 => x"c808b6f8",
   356 => x"1381b72d",
   357 => x"8115558b",
   358 => x"7625ffaa",
   359 => x"38029805",
   360 => x"0d0402fc",
   361 => x"050d7251",
   362 => x"70fd2ead",
   363 => x"3870fd24",
   364 => x"8a3870fc",
   365 => x"2e80c438",
   366 => x"8c830470",
   367 => x"fe2eb138",
   368 => x"70ff2e09",
   369 => x"8106bc38",
   370 => x"b5f80851",
   371 => x"70802eb3",
   372 => x"38ff11b5",
   373 => x"f80c8c83",
   374 => x"04b5f808",
   375 => x"f00570b5",
   376 => x"f80c5170",
   377 => x"80259c38",
   378 => x"800bb5f8",
   379 => x"0c8c8304",
   380 => x"b5f80881",
   381 => x"05b5f80c",
   382 => x"8c8304b5",
   383 => x"f8089005",
   384 => x"b5f80c8a",
   385 => x"872da6c0",
   386 => x"2d028405",
   387 => x"0d0402fc",
   388 => x"050db6f0",
   389 => x"08fb06b6",
   390 => x"f00c7251",
   391 => x"89ce2d02",
   392 => x"84050d04",
   393 => x"02fc050d",
   394 => x"b6f00884",
   395 => x"07b6f00c",
   396 => x"725189ce",
   397 => x"2d028405",
   398 => x"0d0402fc",
   399 => x"050d800b",
   400 => x"b5f80c8a",
   401 => x"872db4c4",
   402 => x"51a7db2d",
   403 => x"b4ac51a7",
   404 => x"eb2d0284",
   405 => x"050d0402",
   406 => x"f8050dbd",
   407 => x"a8088206",
   408 => x"b3dc0b80",
   409 => x"f52d5252",
   410 => x"70802e85",
   411 => x"38718107",
   412 => x"52b3f40b",
   413 => x"80f52d51",
   414 => x"70802e85",
   415 => x"38718407",
   416 => x"52b6f408",
   417 => x"802e8538",
   418 => x"71900752",
   419 => x"71b6c80c",
   420 => x"0288050d",
   421 => x"0402f405",
   422 => x"0d810bb6",
   423 => x"f40c9051",
   424 => x"86922d81",
   425 => x"0bfec40c",
   426 => x"900bfec0",
   427 => x"0c840bfe",
   428 => x"c40c830b",
   429 => x"fecc0ca3",
   430 => x"cb2da5de",
   431 => x"2da3b02d",
   432 => x"a3b02d81",
   433 => x"f72d8151",
   434 => x"84e52da3",
   435 => x"b02da3b0",
   436 => x"2d815184",
   437 => x"e52db1ec",
   438 => x"5185f12d",
   439 => x"84529dc2",
   440 => x"2d8fcc2d",
   441 => x"b6c80880",
   442 => x"2e8638fe",
   443 => x"528df804",
   444 => x"ff125271",
   445 => x"8024e738",
   446 => x"71802e81",
   447 => x"813886c2",
   448 => x"2db28451",
   449 => x"87b42db6",
   450 => x"c808802e",
   451 => x"8f38b3bc",
   452 => x"51a7db2d",
   453 => x"805184e5",
   454 => x"2d8ea604",
   455 => x"b6c80851",
   456 => x"8cba2da5",
   457 => x"ea2da3e3",
   458 => x"2da7f02d",
   459 => x"b6c808bd",
   460 => x"ac08882b",
   461 => x"bdb00807",
   462 => x"fed80c53",
   463 => x"8cd72db6",
   464 => x"c808b6f0",
   465 => x"082ea238",
   466 => x"b6c808b6",
   467 => x"f00cb6c8",
   468 => x"08fec00c",
   469 => x"84527251",
   470 => x"84e52da3",
   471 => x"b02da3b0",
   472 => x"2dff1252",
   473 => x"718025ee",
   474 => x"3872802e",
   475 => x"89388a0b",
   476 => x"fec40c8e",
   477 => x"a604820b",
   478 => x"fec40c8e",
   479 => x"a604b290",
   480 => x"5185f12d",
   481 => x"800bb6c8",
   482 => x"0c028c05",
   483 => x"0d0402e8",
   484 => x"050d7779",
   485 => x"7b585555",
   486 => x"80537276",
   487 => x"25a33874",
   488 => x"70810556",
   489 => x"80f52d74",
   490 => x"70810556",
   491 => x"80f52d52",
   492 => x"5271712e",
   493 => x"86388151",
   494 => x"8fc30481",
   495 => x"13538f9a",
   496 => x"04805170",
   497 => x"b6c80c02",
   498 => x"98050d04",
   499 => x"02d8050d",
   500 => x"800bbcd0",
   501 => x"0cb8c852",
   502 => x"8051a0aa",
   503 => x"2db6c808",
   504 => x"54b6c808",
   505 => x"8c38b2a4",
   506 => x"5185f12d",
   507 => x"735594e7",
   508 => x"04805681",
   509 => x"0bbcf40c",
   510 => x"8853b2b0",
   511 => x"52b8fe51",
   512 => x"8f8e2db6",
   513 => x"c808762e",
   514 => x"09810687",
   515 => x"38b6c808",
   516 => x"bcf40c88",
   517 => x"53b2bc52",
   518 => x"b99a518f",
   519 => x"8e2db6c8",
   520 => x"088738b6",
   521 => x"c808bcf4",
   522 => x"0cbcf408",
   523 => x"802e80f6",
   524 => x"38bc8e0b",
   525 => x"80f52dbc",
   526 => x"8f0b80f5",
   527 => x"2d71982b",
   528 => x"71902b07",
   529 => x"bc900b80",
   530 => x"f52d7088",
   531 => x"2b7207bc",
   532 => x"910b80f5",
   533 => x"2d7107bc",
   534 => x"c60b80f5",
   535 => x"2dbcc70b",
   536 => x"80f52d71",
   537 => x"882b0753",
   538 => x"5f54525a",
   539 => x"56575573",
   540 => x"81abaa2e",
   541 => x"0981068d",
   542 => x"387551a1",
   543 => x"ca2db6c8",
   544 => x"08569192",
   545 => x"047382d4",
   546 => x"d52e8738",
   547 => x"b2c85191",
   548 => x"d304b8c8",
   549 => x"527551a0",
   550 => x"aa2db6c8",
   551 => x"0855b6c8",
   552 => x"08802e83",
   553 => x"c2388853",
   554 => x"b2bc52b9",
   555 => x"9a518f8e",
   556 => x"2db6c808",
   557 => x"8938810b",
   558 => x"bcd00c91",
   559 => x"d9048853",
   560 => x"b2b052b8",
   561 => x"fe518f8e",
   562 => x"2db6c808",
   563 => x"802e8a38",
   564 => x"b2dc5185",
   565 => x"f12d92b3",
   566 => x"04bcc60b",
   567 => x"80f52d54",
   568 => x"7380d52e",
   569 => x"09810680",
   570 => x"ca38bcc7",
   571 => x"0b80f52d",
   572 => x"547381aa",
   573 => x"2e098106",
   574 => x"ba38800b",
   575 => x"b8c80b80",
   576 => x"f52d5654",
   577 => x"7481e92e",
   578 => x"83388154",
   579 => x"7481eb2e",
   580 => x"8c388055",
   581 => x"73752e09",
   582 => x"810682cb",
   583 => x"38b8d30b",
   584 => x"80f52d55",
   585 => x"748d38b8",
   586 => x"d40b80f5",
   587 => x"2d547382",
   588 => x"2e863880",
   589 => x"5594e704",
   590 => x"b8d50b80",
   591 => x"f52d70bc",
   592 => x"c80cff05",
   593 => x"bccc0cb8",
   594 => x"d60b80f5",
   595 => x"2db8d70b",
   596 => x"80f52d58",
   597 => x"76057782",
   598 => x"80290570",
   599 => x"bcd80cb8",
   600 => x"d80b80f5",
   601 => x"2d70bcec",
   602 => x"0cbcd008",
   603 => x"59575876",
   604 => x"802e81a3",
   605 => x"388853b2",
   606 => x"bc52b99a",
   607 => x"518f8e2d",
   608 => x"b6c80881",
   609 => x"e238bcc8",
   610 => x"0870842b",
   611 => x"bcd40c70",
   612 => x"bce80cb8",
   613 => x"ed0b80f5",
   614 => x"2db8ec0b",
   615 => x"80f52d71",
   616 => x"82802905",
   617 => x"b8ee0b80",
   618 => x"f52d7084",
   619 => x"80802912",
   620 => x"b8ef0b80",
   621 => x"f52d7081",
   622 => x"800a2912",
   623 => x"70bcf00c",
   624 => x"bcec0871",
   625 => x"29bcd808",
   626 => x"0570bcdc",
   627 => x"0cb8f50b",
   628 => x"80f52db8",
   629 => x"f40b80f5",
   630 => x"2d718280",
   631 => x"2905b8f6",
   632 => x"0b80f52d",
   633 => x"70848080",
   634 => x"2912b8f7",
   635 => x"0b80f52d",
   636 => x"70982b81",
   637 => x"f00a0672",
   638 => x"0570bce0",
   639 => x"0cfe117e",
   640 => x"297705bc",
   641 => x"e40c5259",
   642 => x"5243545e",
   643 => x"51525952",
   644 => x"5d575957",
   645 => x"94e504b8",
   646 => x"da0b80f5",
   647 => x"2db8d90b",
   648 => x"80f52d71",
   649 => x"82802905",
   650 => x"70bcd40c",
   651 => x"70a02983",
   652 => x"ff057089",
   653 => x"2a70bce8",
   654 => x"0cb8df0b",
   655 => x"80f52db8",
   656 => x"de0b80f5",
   657 => x"2d718280",
   658 => x"290570bc",
   659 => x"f00c7b71",
   660 => x"291e70bc",
   661 => x"e40c7dbc",
   662 => x"e00c7305",
   663 => x"bcdc0c55",
   664 => x"5e515155",
   665 => x"55815574",
   666 => x"b6c80c02",
   667 => x"a8050d04",
   668 => x"02ec050d",
   669 => x"7670872c",
   670 => x"7180ff06",
   671 => x"555654bc",
   672 => x"d0088a38",
   673 => x"73882c74",
   674 => x"81ff0654",
   675 => x"55b8c852",
   676 => x"bcd80815",
   677 => x"51a0aa2d",
   678 => x"b6c80854",
   679 => x"b6c80880",
   680 => x"2eb338bc",
   681 => x"d008802e",
   682 => x"98387284",
   683 => x"29b8c805",
   684 => x"70085253",
   685 => x"a1ca2db6",
   686 => x"c808f00a",
   687 => x"065395d3",
   688 => x"047210b8",
   689 => x"c8057080",
   690 => x"e02d5253",
   691 => x"a1fa2db6",
   692 => x"c8085372",
   693 => x"5473b6c8",
   694 => x"0c029405",
   695 => x"0d0402ec",
   696 => x"050d7670",
   697 => x"842cbce4",
   698 => x"0805718f",
   699 => x"06525553",
   700 => x"728938b8",
   701 => x"c8527351",
   702 => x"a0aa2d72",
   703 => x"a029b8c8",
   704 => x"05548074",
   705 => x"80f52d54",
   706 => x"5572752e",
   707 => x"83388155",
   708 => x"7281e52e",
   709 => x"93387480",
   710 => x"2e8e388b",
   711 => x"1480f52d",
   712 => x"98065372",
   713 => x"802e8338",
   714 => x"805473b6",
   715 => x"c80c0294",
   716 => x"050d0402",
   717 => x"cc050d7e",
   718 => x"605e5a80",
   719 => x"0bbce008",
   720 => x"bce40859",
   721 => x"5c568058",
   722 => x"bcd40878",
   723 => x"2e81ae38",
   724 => x"778f06a0",
   725 => x"17575473",
   726 => x"8f38b8c8",
   727 => x"52765181",
   728 => x"1757a0aa",
   729 => x"2db8c856",
   730 => x"807680f5",
   731 => x"2d565474",
   732 => x"742e8338",
   733 => x"81547481",
   734 => x"e52e80f6",
   735 => x"38817075",
   736 => x"06555c73",
   737 => x"802e80ea",
   738 => x"388b1680",
   739 => x"f52d9806",
   740 => x"597880de",
   741 => x"388b537c",
   742 => x"5275518f",
   743 => x"8e2db6c8",
   744 => x"0880cf38",
   745 => x"9c160851",
   746 => x"a1ca2db6",
   747 => x"c808841b",
   748 => x"0c9a1680",
   749 => x"e02d51a1",
   750 => x"fa2db6c8",
   751 => x"08b6c808",
   752 => x"881c0cb6",
   753 => x"c8085555",
   754 => x"bcd00880",
   755 => x"2e983894",
   756 => x"1680e02d",
   757 => x"51a1fa2d",
   758 => x"b6c80890",
   759 => x"2b83fff0",
   760 => x"0a067016",
   761 => x"51547388",
   762 => x"1b0c787a",
   763 => x"0c7b5498",
   764 => x"b3048118",
   765 => x"58bcd408",
   766 => x"7826fed4",
   767 => x"38bcd008",
   768 => x"802eae38",
   769 => x"7a5194f0",
   770 => x"2db6c808",
   771 => x"b6c80880",
   772 => x"fffffff8",
   773 => x"06555b73",
   774 => x"80ffffff",
   775 => x"f82e9238",
   776 => x"b6c808fe",
   777 => x"05bcc808",
   778 => x"29bcdc08",
   779 => x"055796c6",
   780 => x"04805473",
   781 => x"b6c80c02",
   782 => x"b4050d04",
   783 => x"02f4050d",
   784 => x"74700881",
   785 => x"05710c70",
   786 => x"08bccc08",
   787 => x"06535371",
   788 => x"8e388813",
   789 => x"085194f0",
   790 => x"2db6c808",
   791 => x"88140c81",
   792 => x"0bb6c80c",
   793 => x"028c050d",
   794 => x"0402f005",
   795 => x"0d758811",
   796 => x"08fe05bc",
   797 => x"c80829bc",
   798 => x"dc081172",
   799 => x"08bccc08",
   800 => x"06057955",
   801 => x"535454a0",
   802 => x"aa2d0290",
   803 => x"050d0402",
   804 => x"f0050d75",
   805 => x"881108fe",
   806 => x"05bcc808",
   807 => x"29bcdc08",
   808 => x"117208bc",
   809 => x"cc080605",
   810 => x"79555354",
   811 => x"549eea2d",
   812 => x"0290050d",
   813 => x"0402f405",
   814 => x"0dd45281",
   815 => x"ff720c71",
   816 => x"085381ff",
   817 => x"720c7288",
   818 => x"2b83fe80",
   819 => x"06720870",
   820 => x"81ff0651",
   821 => x"525381ff",
   822 => x"720c7271",
   823 => x"07882b72",
   824 => x"087081ff",
   825 => x"06515253",
   826 => x"81ff720c",
   827 => x"72710788",
   828 => x"2b720870",
   829 => x"81ff0672",
   830 => x"07b6c80c",
   831 => x"5253028c",
   832 => x"050d0402",
   833 => x"f4050d74",
   834 => x"767181ff",
   835 => x"06d40c53",
   836 => x"53bcf808",
   837 => x"85387189",
   838 => x"2b527198",
   839 => x"2ad40c71",
   840 => x"902a7081",
   841 => x"ff06d40c",
   842 => x"5171882a",
   843 => x"7081ff06",
   844 => x"d40c5171",
   845 => x"81ff06d4",
   846 => x"0c72902a",
   847 => x"7081ff06",
   848 => x"d40c51d4",
   849 => x"087081ff",
   850 => x"06515182",
   851 => x"b8bf5270",
   852 => x"81ff2e09",
   853 => x"81069438",
   854 => x"81ff0bd4",
   855 => x"0cd40870",
   856 => x"81ff06ff",
   857 => x"14545151",
   858 => x"71e53870",
   859 => x"b6c80c02",
   860 => x"8c050d04",
   861 => x"02fc050d",
   862 => x"81c75181",
   863 => x"ff0bd40c",
   864 => x"ff115170",
   865 => x"8025f438",
   866 => x"0284050d",
   867 => x"0402f005",
   868 => x"0d9af42d",
   869 => x"8fcf5380",
   870 => x"5287fc80",
   871 => x"f7519a83",
   872 => x"2db6c808",
   873 => x"54b6c808",
   874 => x"812e0981",
   875 => x"06a33881",
   876 => x"ff0bd40c",
   877 => x"820a5284",
   878 => x"9c80e951",
   879 => x"9a832db6",
   880 => x"c8088b38",
   881 => x"81ff0bd4",
   882 => x"0c73539b",
   883 => x"d7049af4",
   884 => x"2dff1353",
   885 => x"72c13872",
   886 => x"b6c80c02",
   887 => x"90050d04",
   888 => x"02f4050d",
   889 => x"81ff0bd4",
   890 => x"0c935380",
   891 => x"5287fc80",
   892 => x"c1519a83",
   893 => x"2db6c808",
   894 => x"8b3881ff",
   895 => x"0bd40c81",
   896 => x"539c8d04",
   897 => x"9af42dff",
   898 => x"135372df",
   899 => x"3872b6c8",
   900 => x"0c028c05",
   901 => x"0d0402f0",
   902 => x"050d9af4",
   903 => x"2d83aa52",
   904 => x"849c80c8",
   905 => x"519a832d",
   906 => x"b6c80881",
   907 => x"2e098106",
   908 => x"923899b5",
   909 => x"2db6c808",
   910 => x"83ffff06",
   911 => x"537283aa",
   912 => x"2e97389b",
   913 => x"e02d9cd4",
   914 => x"0481549d",
   915 => x"b904b2e8",
   916 => x"5185f12d",
   917 => x"80549db9",
   918 => x"0481ff0b",
   919 => x"d40cb153",
   920 => x"9b8d2db6",
   921 => x"c808802e",
   922 => x"80c03880",
   923 => x"5287fc80",
   924 => x"fa519a83",
   925 => x"2db6c808",
   926 => x"b13881ff",
   927 => x"0bd40cd4",
   928 => x"085381ff",
   929 => x"0bd40c81",
   930 => x"ff0bd40c",
   931 => x"81ff0bd4",
   932 => x"0c81ff0b",
   933 => x"d40c7286",
   934 => x"2a708106",
   935 => x"b6c80856",
   936 => x"51537280",
   937 => x"2e93389c",
   938 => x"c9047282",
   939 => x"2eff9f38",
   940 => x"ff135372",
   941 => x"ffaa3872",
   942 => x"5473b6c8",
   943 => x"0c029005",
   944 => x"0d0402f0",
   945 => x"050d810b",
   946 => x"bcf80c84",
   947 => x"54d00870",
   948 => x"8f2a7081",
   949 => x"06515153",
   950 => x"72f33872",
   951 => x"d00c9af4",
   952 => x"2db2f851",
   953 => x"85f12dd0",
   954 => x"08708f2a",
   955 => x"70810651",
   956 => x"515372f3",
   957 => x"38810bd0",
   958 => x"0cb15380",
   959 => x"5284d480",
   960 => x"c0519a83",
   961 => x"2db6c808",
   962 => x"812ea138",
   963 => x"72822e09",
   964 => x"81068c38",
   965 => x"b3845185",
   966 => x"f12d8053",
   967 => x"9ee104ff",
   968 => x"135372d7",
   969 => x"38ff1454",
   970 => x"73ffa238",
   971 => x"9c962db6",
   972 => x"c808bcf8",
   973 => x"0cb6c808",
   974 => x"8b388152",
   975 => x"87fc80d0",
   976 => x"519a832d",
   977 => x"81ff0bd4",
   978 => x"0cd00870",
   979 => x"8f2a7081",
   980 => x"06515153",
   981 => x"72f33872",
   982 => x"d00c81ff",
   983 => x"0bd40c81",
   984 => x"5372b6c8",
   985 => x"0c029005",
   986 => x"0d0402e8",
   987 => x"050d7856",
   988 => x"81ff0bd4",
   989 => x"0cd00870",
   990 => x"8f2a7081",
   991 => x"06515153",
   992 => x"72f33882",
   993 => x"810bd00c",
   994 => x"81ff0bd4",
   995 => x"0c775287",
   996 => x"fc80d851",
   997 => x"9a832db6",
   998 => x"c808802e",
   999 => x"8c38b39c",
  1000 => x"5185f12d",
  1001 => x"8153a0a1",
  1002 => x"0481ff0b",
  1003 => x"d40c81fe",
  1004 => x"0bd40c80",
  1005 => x"ff557570",
  1006 => x"84055708",
  1007 => x"70982ad4",
  1008 => x"0c70902c",
  1009 => x"7081ff06",
  1010 => x"d40c5470",
  1011 => x"882c7081",
  1012 => x"ff06d40c",
  1013 => x"547081ff",
  1014 => x"06d40c54",
  1015 => x"ff155574",
  1016 => x"8025d338",
  1017 => x"81ff0bd4",
  1018 => x"0c81ff0b",
  1019 => x"d40c81ff",
  1020 => x"0bd40c86",
  1021 => x"8da05481",
  1022 => x"ff0bd40c",
  1023 => x"d40881ff",
  1024 => x"06557487",
  1025 => x"38ff1454",
  1026 => x"73ed3881",
  1027 => x"ff0bd40c",
  1028 => x"d008708f",
  1029 => x"2a708106",
  1030 => x"51515372",
  1031 => x"f33872d0",
  1032 => x"0c72b6c8",
  1033 => x"0c029805",
  1034 => x"0d0402e8",
  1035 => x"050d7855",
  1036 => x"805681ff",
  1037 => x"0bd40cd0",
  1038 => x"08708f2a",
  1039 => x"70810651",
  1040 => x"515372f3",
  1041 => x"3882810b",
  1042 => x"d00c81ff",
  1043 => x"0bd40c77",
  1044 => x"5287fc80",
  1045 => x"d1519a83",
  1046 => x"2d80dbc6",
  1047 => x"df54b6c8",
  1048 => x"08802e8a",
  1049 => x"38b1d451",
  1050 => x"85f12da1",
  1051 => x"c10481ff",
  1052 => x"0bd40cd4",
  1053 => x"087081ff",
  1054 => x"06515372",
  1055 => x"81fe2e09",
  1056 => x"81069d38",
  1057 => x"80ff5399",
  1058 => x"b52db6c8",
  1059 => x"08757084",
  1060 => x"05570cff",
  1061 => x"13537280",
  1062 => x"25ed3881",
  1063 => x"56a1a604",
  1064 => x"ff145473",
  1065 => x"c93881ff",
  1066 => x"0bd40c81",
  1067 => x"ff0bd40c",
  1068 => x"d008708f",
  1069 => x"2a708106",
  1070 => x"51515372",
  1071 => x"f33872d0",
  1072 => x"0c75b6c8",
  1073 => x"0c029805",
  1074 => x"0d0402f4",
  1075 => x"050d7470",
  1076 => x"882a83fe",
  1077 => x"80067072",
  1078 => x"982a0772",
  1079 => x"882b87fc",
  1080 => x"80800673",
  1081 => x"982b81f0",
  1082 => x"0a067173",
  1083 => x"0707b6c8",
  1084 => x"0c565153",
  1085 => x"51028c05",
  1086 => x"0d0402f8",
  1087 => x"050d028e",
  1088 => x"0580f52d",
  1089 => x"74882b07",
  1090 => x"7083ffff",
  1091 => x"06b6c80c",
  1092 => x"51028805",
  1093 => x"0d0402fc",
  1094 => x"050d7251",
  1095 => x"80710c80",
  1096 => x"0b84120c",
  1097 => x"0284050d",
  1098 => x"0402f005",
  1099 => x"0d757008",
  1100 => x"84120853",
  1101 => x"5353ff54",
  1102 => x"71712ea8",
  1103 => x"38a5e42d",
  1104 => x"84130870",
  1105 => x"84291488",
  1106 => x"11700870",
  1107 => x"81ff0684",
  1108 => x"18088111",
  1109 => x"8706841a",
  1110 => x"0c535155",
  1111 => x"515151a5",
  1112 => x"de2d7154",
  1113 => x"73b6c80c",
  1114 => x"0290050d",
  1115 => x"0402f805",
  1116 => x"0da5e42d",
  1117 => x"e008708b",
  1118 => x"2a708106",
  1119 => x"51525270",
  1120 => x"802e9d38",
  1121 => x"bcfc0870",
  1122 => x"8429bd84",
  1123 => x"057381ff",
  1124 => x"06710c51",
  1125 => x"51bcfc08",
  1126 => x"81118706",
  1127 => x"bcfc0c51",
  1128 => x"800bbda4",
  1129 => x"0ca5d72d",
  1130 => x"a5de2d02",
  1131 => x"88050d04",
  1132 => x"02fc050d",
  1133 => x"a5e42d81",
  1134 => x"0bbda40c",
  1135 => x"a5de2dbd",
  1136 => x"a4085170",
  1137 => x"fa380284",
  1138 => x"050d0402",
  1139 => x"fc050dbc",
  1140 => x"fc51a296",
  1141 => x"2da2ed51",
  1142 => x"a5d32da4",
  1143 => x"fd2d0284",
  1144 => x"050d0402",
  1145 => x"f4050da4",
  1146 => x"e504b6c8",
  1147 => x"0881f02e",
  1148 => x"09810689",
  1149 => x"38810bb6",
  1150 => x"bc0ca4e5",
  1151 => x"04b6c808",
  1152 => x"81e02e09",
  1153 => x"81068938",
  1154 => x"810bb6c0",
  1155 => x"0ca4e504",
  1156 => x"b6c80852",
  1157 => x"b6c00880",
  1158 => x"2e8838b6",
  1159 => x"c8088180",
  1160 => x"05527184",
  1161 => x"2c728f06",
  1162 => x"5353b6bc",
  1163 => x"08802e99",
  1164 => x"38728429",
  1165 => x"b5fc0572",
  1166 => x"1381712b",
  1167 => x"70097308",
  1168 => x"06730c51",
  1169 => x"5353a4db",
  1170 => x"04728429",
  1171 => x"b5fc0572",
  1172 => x"1383712b",
  1173 => x"72080772",
  1174 => x"0c535380",
  1175 => x"0bb6c00c",
  1176 => x"800bb6bc",
  1177 => x"0cbcfc51",
  1178 => x"a2a92db6",
  1179 => x"c808ff24",
  1180 => x"fef83880",
  1181 => x"0bb6c80c",
  1182 => x"028c050d",
  1183 => x"0402f805",
  1184 => x"0db5fc52",
  1185 => x"8f518072",
  1186 => x"70840554",
  1187 => x"0cff1151",
  1188 => x"708025f2",
  1189 => x"38028805",
  1190 => x"0d0402f0",
  1191 => x"050d7551",
  1192 => x"a5e42d70",
  1193 => x"822cfc06",
  1194 => x"b5fc1172",
  1195 => x"109e0671",
  1196 => x"0870722a",
  1197 => x"70830682",
  1198 => x"742b7009",
  1199 => x"7406760c",
  1200 => x"54515657",
  1201 => x"535153a5",
  1202 => x"de2d71b6",
  1203 => x"c80c0290",
  1204 => x"050d0471",
  1205 => x"980c04ff",
  1206 => x"b008b6c8",
  1207 => x"0c04810b",
  1208 => x"ffb00c04",
  1209 => x"800bffb0",
  1210 => x"0c0402fc",
  1211 => x"050d810b",
  1212 => x"b6c40c81",
  1213 => x"5184e52d",
  1214 => x"0284050d",
  1215 => x"0402fc05",
  1216 => x"0d800bb6",
  1217 => x"c40c8051",
  1218 => x"84e52d02",
  1219 => x"84050d04",
  1220 => x"02ec050d",
  1221 => x"76548052",
  1222 => x"870b8815",
  1223 => x"80f52d56",
  1224 => x"53747224",
  1225 => x"8338a053",
  1226 => x"725182ee",
  1227 => x"2d81128b",
  1228 => x"1580f52d",
  1229 => x"54527272",
  1230 => x"25de3802",
  1231 => x"94050d04",
  1232 => x"02f0050d",
  1233 => x"bdb40854",
  1234 => x"81f72d80",
  1235 => x"0bbdb80c",
  1236 => x"7308802e",
  1237 => x"81803882",
  1238 => x"0bb6dc0c",
  1239 => x"bdb8088f",
  1240 => x"06b6d80c",
  1241 => x"73085271",
  1242 => x"832e9638",
  1243 => x"71832689",
  1244 => x"3871812e",
  1245 => x"af38a7c1",
  1246 => x"0471852e",
  1247 => x"9f38a7c1",
  1248 => x"04881480",
  1249 => x"f52d8415",
  1250 => x"08b3ac53",
  1251 => x"545285f1",
  1252 => x"2d718429",
  1253 => x"13700852",
  1254 => x"52a7c504",
  1255 => x"7351a690",
  1256 => x"2da7c104",
  1257 => x"bda80888",
  1258 => x"15082c70",
  1259 => x"81065152",
  1260 => x"71802e87",
  1261 => x"38b3b051",
  1262 => x"a7be04b3",
  1263 => x"b45185f1",
  1264 => x"2d841408",
  1265 => x"5185f12d",
  1266 => x"bdb80881",
  1267 => x"05bdb80c",
  1268 => x"8c1454a6",
  1269 => x"d0040290",
  1270 => x"050d0471",
  1271 => x"bdb40ca6",
  1272 => x"c02dbdb8",
  1273 => x"08ff05bd",
  1274 => x"bc0c0471",
  1275 => x"bdc00c04",
  1276 => x"02e8050d",
  1277 => x"bdb408bd",
  1278 => x"c0085755",
  1279 => x"80f851a5",
  1280 => x"9a2db6c8",
  1281 => x"08812a70",
  1282 => x"81065152",
  1283 => x"719b3887",
  1284 => x"51a59a2d",
  1285 => x"b6c80881",
  1286 => x"2a708106",
  1287 => x"51527180",
  1288 => x"2eb138a8",
  1289 => x"a904a3e3",
  1290 => x"2d8751a5",
  1291 => x"9a2db6c8",
  1292 => x"08f438a8",
  1293 => x"b904a3e3",
  1294 => x"2d80f851",
  1295 => x"a59a2db6",
  1296 => x"c808f338",
  1297 => x"b6c40881",
  1298 => x"3270b6c4",
  1299 => x"0c705252",
  1300 => x"84e52d80",
  1301 => x"0bbdac0c",
  1302 => x"800bbdb0",
  1303 => x"0cb6c408",
  1304 => x"82dd3880",
  1305 => x"da51a59a",
  1306 => x"2db6c808",
  1307 => x"802e8a38",
  1308 => x"bdac0881",
  1309 => x"8007bdac",
  1310 => x"0c80d951",
  1311 => x"a59a2db6",
  1312 => x"c808802e",
  1313 => x"8a38bdac",
  1314 => x"0880c007",
  1315 => x"bdac0c81",
  1316 => x"9451a59a",
  1317 => x"2db6c808",
  1318 => x"802e8938",
  1319 => x"bdac0890",
  1320 => x"07bdac0c",
  1321 => x"819151a5",
  1322 => x"9a2db6c8",
  1323 => x"08802e89",
  1324 => x"38bdac08",
  1325 => x"a007bdac",
  1326 => x"0c81f551",
  1327 => x"a59a2db6",
  1328 => x"c808802e",
  1329 => x"8938bdac",
  1330 => x"088107bd",
  1331 => x"ac0c81f2",
  1332 => x"51a59a2d",
  1333 => x"b6c80880",
  1334 => x"2e8938bd",
  1335 => x"ac088207",
  1336 => x"bdac0c81",
  1337 => x"eb51a59a",
  1338 => x"2db6c808",
  1339 => x"802e8938",
  1340 => x"bdac0884",
  1341 => x"07bdac0c",
  1342 => x"81f451a5",
  1343 => x"9a2db6c8",
  1344 => x"08802e89",
  1345 => x"38bdac08",
  1346 => x"8807bdac",
  1347 => x"0c80d851",
  1348 => x"a59a2db6",
  1349 => x"c808802e",
  1350 => x"8a38bdb0",
  1351 => x"08818007",
  1352 => x"bdb00c92",
  1353 => x"51a59a2d",
  1354 => x"b6c80880",
  1355 => x"2e8a38bd",
  1356 => x"b00880c0",
  1357 => x"07bdb00c",
  1358 => x"9451a59a",
  1359 => x"2db6c808",
  1360 => x"802e8938",
  1361 => x"bdb00890",
  1362 => x"07bdb00c",
  1363 => x"9151a59a",
  1364 => x"2db6c808",
  1365 => x"802e8938",
  1366 => x"bdb008a0",
  1367 => x"07bdb00c",
  1368 => x"9d51a59a",
  1369 => x"2db6c808",
  1370 => x"802e8938",
  1371 => x"bdb00881",
  1372 => x"07bdb00c",
  1373 => x"9b51a59a",
  1374 => x"2db6c808",
  1375 => x"802e8938",
  1376 => x"bdb00882",
  1377 => x"07bdb00c",
  1378 => x"9c51a59a",
  1379 => x"2db6c808",
  1380 => x"802e8938",
  1381 => x"bdb00884",
  1382 => x"07bdb00c",
  1383 => x"a351a59a",
  1384 => x"2db6c808",
  1385 => x"802e8938",
  1386 => x"bdb00888",
  1387 => x"07bdb00c",
  1388 => x"81fd51a5",
  1389 => x"9a2d81fa",
  1390 => x"51a59a2d",
  1391 => x"b0a40481",
  1392 => x"f551a59a",
  1393 => x"2db6c808",
  1394 => x"812a7081",
  1395 => x"06515271",
  1396 => x"802eaf38",
  1397 => x"bdbc0852",
  1398 => x"71802e89",
  1399 => x"38ff12bd",
  1400 => x"bc0cac82",
  1401 => x"04bdb808",
  1402 => x"10bdb808",
  1403 => x"05708429",
  1404 => x"16515288",
  1405 => x"1208802e",
  1406 => x"8938ff51",
  1407 => x"88120852",
  1408 => x"712d81f2",
  1409 => x"51a59a2d",
  1410 => x"b6c80881",
  1411 => x"2a708106",
  1412 => x"51527180",
  1413 => x"2eb138bd",
  1414 => x"b808ff11",
  1415 => x"bdbc0856",
  1416 => x"53537372",
  1417 => x"25893881",
  1418 => x"14bdbc0c",
  1419 => x"acc70472",
  1420 => x"10137084",
  1421 => x"29165152",
  1422 => x"88120880",
  1423 => x"2e8938fe",
  1424 => x"51881208",
  1425 => x"52712d81",
  1426 => x"fd51a59a",
  1427 => x"2db6c808",
  1428 => x"812a7081",
  1429 => x"06515271",
  1430 => x"802e8638",
  1431 => x"800bbdbc",
  1432 => x"0c81fa51",
  1433 => x"a59a2db6",
  1434 => x"c808812a",
  1435 => x"70810651",
  1436 => x"5271802e",
  1437 => x"8938bdb8",
  1438 => x"08ff05bd",
  1439 => x"bc0cbdbc",
  1440 => x"08705354",
  1441 => x"73802e8a",
  1442 => x"388c15ff",
  1443 => x"155555ad",
  1444 => x"8404820b",
  1445 => x"b6dc0c71",
  1446 => x"8f06b6d8",
  1447 => x"0c81eb51",
  1448 => x"a59a2db6",
  1449 => x"c808812a",
  1450 => x"70810651",
  1451 => x"5271802e",
  1452 => x"ad387408",
  1453 => x"852e0981",
  1454 => x"06a43888",
  1455 => x"1580f52d",
  1456 => x"ff055271",
  1457 => x"881681b7",
  1458 => x"2d71982b",
  1459 => x"52718025",
  1460 => x"8838800b",
  1461 => x"881681b7",
  1462 => x"2d7451a6",
  1463 => x"902d81f4",
  1464 => x"51a59a2d",
  1465 => x"b6c80881",
  1466 => x"2a708106",
  1467 => x"51527180",
  1468 => x"2eb33874",
  1469 => x"08852e09",
  1470 => x"8106aa38",
  1471 => x"881580f5",
  1472 => x"2d810552",
  1473 => x"71881681",
  1474 => x"b72d7181",
  1475 => x"ff068b16",
  1476 => x"80f52d54",
  1477 => x"52727227",
  1478 => x"87387288",
  1479 => x"1681b72d",
  1480 => x"7451a690",
  1481 => x"2d80da51",
  1482 => x"a59a2db6",
  1483 => x"c808812a",
  1484 => x"70810651",
  1485 => x"5271802e",
  1486 => x"81a638bd",
  1487 => x"b408bdbc",
  1488 => x"08555373",
  1489 => x"802e8a38",
  1490 => x"8c13ff15",
  1491 => x"5553aec3",
  1492 => x"04720852",
  1493 => x"71822ea6",
  1494 => x"38718226",
  1495 => x"89387181",
  1496 => x"2ea938af",
  1497 => x"e0047183",
  1498 => x"2eb13871",
  1499 => x"842e0981",
  1500 => x"0680ed38",
  1501 => x"88130851",
  1502 => x"a7db2daf",
  1503 => x"e004bdbc",
  1504 => x"08518813",
  1505 => x"0852712d",
  1506 => x"afe00481",
  1507 => x"0b881408",
  1508 => x"2bbda808",
  1509 => x"32bda80c",
  1510 => x"afb60488",
  1511 => x"1380f52d",
  1512 => x"81058b14",
  1513 => x"80f52d53",
  1514 => x"54717424",
  1515 => x"83388054",
  1516 => x"73881481",
  1517 => x"b72da6c0",
  1518 => x"2dafe004",
  1519 => x"7508802e",
  1520 => x"a2387508",
  1521 => x"51a59a2d",
  1522 => x"b6c80881",
  1523 => x"06527180",
  1524 => x"2e8b38bd",
  1525 => x"bc085184",
  1526 => x"16085271",
  1527 => x"2d881656",
  1528 => x"75da3880",
  1529 => x"54800bb6",
  1530 => x"dc0c738f",
  1531 => x"06b6d80c",
  1532 => x"a05273bd",
  1533 => x"bc082e09",
  1534 => x"81069838",
  1535 => x"bdb808ff",
  1536 => x"05743270",
  1537 => x"09810570",
  1538 => x"72079f2a",
  1539 => x"91713151",
  1540 => x"51535371",
  1541 => x"5182ee2d",
  1542 => x"8114548e",
  1543 => x"7425c638",
  1544 => x"b6c40852",
  1545 => x"71b6c80c",
  1546 => x"0298050d",
  1547 => x"04000000",
  1548 => x"00ffffff",
  1549 => x"ff00ffff",
  1550 => x"ffff00ff",
  1551 => x"ffffff00",
  1552 => x"52657365",
  1553 => x"74000000",
  1554 => x"53617665",
  1555 => x"20736574",
  1556 => x"74696e67",
  1557 => x"73000000",
  1558 => x"5363616e",
  1559 => x"6c696e65",
  1560 => x"73000000",
  1561 => x"4c6f6164",
  1562 => x"20524f4d",
  1563 => x"20100000",
  1564 => x"45786974",
  1565 => x"00000000",
  1566 => x"50432045",
  1567 => x"6e67696e",
  1568 => x"65206d6f",
  1569 => x"64650000",
  1570 => x"54757262",
  1571 => x"6f677261",
  1572 => x"66782031",
  1573 => x"36206d6f",
  1574 => x"64650000",
  1575 => x"56474120",
  1576 => x"2d203331",
  1577 => x"4b487a2c",
  1578 => x"20363048",
  1579 => x"7a000000",
  1580 => x"5456202d",
  1581 => x"20343830",
  1582 => x"692c2036",
  1583 => x"30487a00",
  1584 => x"4261636b",
  1585 => x"00000000",
  1586 => x"46504741",
  1587 => x"50434520",
  1588 => x"43464700",
  1589 => x"52656164",
  1590 => x"20666169",
  1591 => x"6c65640a",
  1592 => x"00000000",
  1593 => x"4661696c",
  1594 => x"65640a00",
  1595 => x"496e6974",
  1596 => x"69616c69",
  1597 => x"7a696e67",
  1598 => x"20534420",
  1599 => x"63617264",
  1600 => x"0a000000",
  1601 => x"424f4f54",
  1602 => x"20202020",
  1603 => x"50434500",
  1604 => x"43617264",
  1605 => x"20696e69",
  1606 => x"74206661",
  1607 => x"696c6564",
  1608 => x"0a000000",
  1609 => x"4d425220",
  1610 => x"6661696c",
  1611 => x"0a000000",
  1612 => x"46415431",
  1613 => x"36202020",
  1614 => x"00000000",
  1615 => x"46415433",
  1616 => x"32202020",
  1617 => x"00000000",
  1618 => x"4e6f2070",
  1619 => x"61727469",
  1620 => x"74696f6e",
  1621 => x"20736967",
  1622 => x"0a000000",
  1623 => x"42616420",
  1624 => x"70617274",
  1625 => x"0a000000",
  1626 => x"53444843",
  1627 => x"20657272",
  1628 => x"6f72210a",
  1629 => x"00000000",
  1630 => x"53442069",
  1631 => x"6e69742e",
  1632 => x"2e2e0a00",
  1633 => x"53442063",
  1634 => x"61726420",
  1635 => x"72657365",
  1636 => x"74206661",
  1637 => x"696c6564",
  1638 => x"210a0000",
  1639 => x"57726974",
  1640 => x"65206661",
  1641 => x"696c6564",
  1642 => x"0a000000",
  1643 => x"16200000",
  1644 => x"14200000",
  1645 => x"15200000",
  1646 => x"00000002",
  1647 => x"00000002",
  1648 => x"00001840",
  1649 => x"000004b9",
  1650 => x"00000002",
  1651 => x"00001848",
  1652 => x"00000377",
  1653 => x"00000003",
  1654 => x"00001a24",
  1655 => x"00000002",
  1656 => x"00000001",
  1657 => x"00001858",
  1658 => x"00000002",
  1659 => x"00000003",
  1660 => x"00001a1c",
  1661 => x"00000002",
  1662 => x"00000002",
  1663 => x"00001864",
  1664 => x"0000063a",
  1665 => x"00000002",
  1666 => x"00001870",
  1667 => x"000012fd",
  1668 => x"00000000",
  1669 => x"00000000",
  1670 => x"00000000",
  1671 => x"00001878",
  1672 => x"00001888",
  1673 => x"0000189c",
  1674 => x"000018b0",
  1675 => x"0000004d",
  1676 => x"0000060e",
  1677 => x"0000002c",
  1678 => x"00000624",
  1679 => x"00000000",
  1680 => x"00000000",
  1681 => x"00000002",
  1682 => x"00001b78",
  1683 => x"000004ce",
  1684 => x"00000002",
  1685 => x"00001b88",
  1686 => x"000004ce",
  1687 => x"00000002",
  1688 => x"00001b98",
  1689 => x"000004ce",
  1690 => x"00000002",
  1691 => x"00001ba8",
  1692 => x"000004ce",
  1693 => x"00000002",
  1694 => x"00001bb8",
  1695 => x"000004ce",
  1696 => x"00000002",
  1697 => x"00001bc8",
  1698 => x"000004ce",
  1699 => x"00000002",
  1700 => x"00001bd8",
  1701 => x"000004ce",
  1702 => x"00000002",
  1703 => x"00001be8",
  1704 => x"000004ce",
  1705 => x"00000002",
  1706 => x"00001bf8",
  1707 => x"000004ce",
  1708 => x"00000002",
  1709 => x"00001c08",
  1710 => x"000004ce",
  1711 => x"00000002",
  1712 => x"00001c18",
  1713 => x"000004ce",
  1714 => x"00000002",
  1715 => x"00001c28",
  1716 => x"000004ce",
  1717 => x"00000002",
  1718 => x"00001c38",
  1719 => x"000004ce",
  1720 => x"00000004",
  1721 => x"000018c0",
  1722 => x"000019bc",
  1723 => x"00000000",
  1724 => x"00000000",
  1725 => x"000005a2",
  1726 => x"00000000",
  1727 => x"00000000",
  1728 => x"00000000",
  1729 => x"00000000",
  1730 => x"00000000",
  1731 => x"00000000",
  1732 => x"00000000",
  1733 => x"00000000",
  1734 => x"00000000",
  1735 => x"00000000",
  1736 => x"00000000",
  1737 => x"00000000",
  1738 => x"00000000",
  1739 => x"00000000",
  1740 => x"00000000",
  1741 => x"00000000",
  1742 => x"00000000",
  1743 => x"00000000",
  1744 => x"00000000",
  1745 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

