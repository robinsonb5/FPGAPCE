-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bbd",
     9 => x"ec080b0b",
    10 => x"0bbdf008",
    11 => x"0b0b0bbd",
    12 => x"f4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bdf40c0b",
    16 => x"0b0bbdf0",
    17 => x"0c0b0b0b",
    18 => x"bdec0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb7d8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bdec7080",
    57 => x"c8ac278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"518fce04",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbdfc0c",
    65 => x"9f0bbe80",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"be8008ff",
    69 => x"05be800c",
    70 => x"be800880",
    71 => x"25eb38bd",
    72 => x"fc08ff05",
    73 => x"bdfc0cbd",
    74 => x"fc088025",
    75 => x"d7380284",
    76 => x"050d0402",
    77 => x"f0050df8",
    78 => x"8053f8a0",
    79 => x"5483bf52",
    80 => x"73708105",
    81 => x"55335170",
    82 => x"73708105",
    83 => x"5534ff12",
    84 => x"52718025",
    85 => x"eb38fbc0",
    86 => x"539f52a0",
    87 => x"73708105",
    88 => x"5534ff12",
    89 => x"52718025",
    90 => x"f2380290",
    91 => x"050d0402",
    92 => x"f4050d74",
    93 => x"538e0bbd",
    94 => x"fc08258f",
    95 => x"3882b32d",
    96 => x"bdfc08ff",
    97 => x"05bdfc0c",
    98 => x"82f504bd",
    99 => x"fc08be80",
   100 => x"08535172",
   101 => x"8a2e0981",
   102 => x"06b73871",
   103 => x"51719f24",
   104 => x"a038bdfc",
   105 => x"08a02911",
   106 => x"f8801151",
   107 => x"51a07134",
   108 => x"be800881",
   109 => x"05be800c",
   110 => x"be800851",
   111 => x"9f7125e2",
   112 => x"38800bbe",
   113 => x"800cbdfc",
   114 => x"088105bd",
   115 => x"fc0c83e5",
   116 => x"0470a029",
   117 => x"12f88011",
   118 => x"51517271",
   119 => x"34be8008",
   120 => x"8105be80",
   121 => x"0cbe8008",
   122 => x"a02e0981",
   123 => x"068e3880",
   124 => x"0bbe800c",
   125 => x"bdfc0881",
   126 => x"05bdfc0c",
   127 => x"028c050d",
   128 => x"0402e805",
   129 => x"0d777956",
   130 => x"56880bfc",
   131 => x"1677712c",
   132 => x"8f065452",
   133 => x"54805372",
   134 => x"72259538",
   135 => x"7153fbe0",
   136 => x"14518771",
   137 => x"348114ff",
   138 => x"14545472",
   139 => x"f1387153",
   140 => x"f9157671",
   141 => x"2c870653",
   142 => x"5171802e",
   143 => x"8b38fbe0",
   144 => x"14517171",
   145 => x"34811454",
   146 => x"728e2495",
   147 => x"388f7331",
   148 => x"53fbe014",
   149 => x"51a07134",
   150 => x"8114ff14",
   151 => x"545472f1",
   152 => x"38029805",
   153 => x"0d0402ec",
   154 => x"050d800b",
   155 => x"be840cf6",
   156 => x"8c08f690",
   157 => x"0871882c",
   158 => x"565481ff",
   159 => x"06527372",
   160 => x"25883871",
   161 => x"54820bbe",
   162 => x"840c7288",
   163 => x"2c7381ff",
   164 => x"06545574",
   165 => x"73258b38",
   166 => x"72be8408",
   167 => x"8407be84",
   168 => x"0c557384",
   169 => x"2b87e871",
   170 => x"25837131",
   171 => x"700b0b0b",
   172 => x"bad80c81",
   173 => x"712bf688",
   174 => x"0cfea413",
   175 => x"ff122c78",
   176 => x"8829ff94",
   177 => x"0570812c",
   178 => x"be840852",
   179 => x"58525551",
   180 => x"52547680",
   181 => x"2e853870",
   182 => x"81075170",
   183 => x"f6940c71",
   184 => x"098105f6",
   185 => x"800c7209",
   186 => x"8105f684",
   187 => x"0c029405",
   188 => x"0d0402f4",
   189 => x"050d7453",
   190 => x"72708105",
   191 => x"5480f52d",
   192 => x"5271802e",
   193 => x"89387151",
   194 => x"82ef2d85",
   195 => x"f804028c",
   196 => x"050d0402",
   197 => x"f4050d74",
   198 => x"70820680",
   199 => x"c8900cba",
   200 => x"f4718106",
   201 => x"54545171",
   202 => x"881481b7",
   203 => x"2d70822a",
   204 => x"70810651",
   205 => x"5170a014",
   206 => x"81b72d70",
   207 => x"bdec0c02",
   208 => x"8c050d04",
   209 => x"02f8050d",
   210 => x"b8f052be",
   211 => x"88519caf",
   212 => x"2dbdec08",
   213 => x"802ea138",
   214 => x"80c1a452",
   215 => x"be88519e",
   216 => x"f02d80c1",
   217 => x"a408be94",
   218 => x"0c80c1a4",
   219 => x"08fec00c",
   220 => x"80c1a408",
   221 => x"5186932d",
   222 => x"0288050d",
   223 => x"0402f005",
   224 => x"0d805192",
   225 => x"872db8f0",
   226 => x"52be8851",
   227 => x"9caf2dbd",
   228 => x"ec08802e",
   229 => x"a838be94",
   230 => x"0880c1a4",
   231 => x"0c80c1a8",
   232 => x"5480fd53",
   233 => x"80747084",
   234 => x"05560cff",
   235 => x"13537280",
   236 => x"25f23880",
   237 => x"c1a452be",
   238 => x"88519f99",
   239 => x"2d029005",
   240 => x"0d0402d4",
   241 => x"050dbe94",
   242 => x"08fec00c",
   243 => x"810bfec4",
   244 => x"0c840bfe",
   245 => x"c40c7c52",
   246 => x"be88519c",
   247 => x"af2dbdec",
   248 => x"0853bdec",
   249 => x"08802e81",
   250 => x"ce38be8c",
   251 => x"0856800b",
   252 => x"ff175859",
   253 => x"76792e8b",
   254 => x"38811977",
   255 => x"812a5859",
   256 => x"76f738f7",
   257 => x"19769fff",
   258 => x"06545972",
   259 => x"802e8b38",
   260 => x"fc8016be",
   261 => x"8852569e",
   262 => x"c22d75b0",
   263 => x"80802e09",
   264 => x"81068938",
   265 => x"820bfedc",
   266 => x"0c88c304",
   267 => x"75988080",
   268 => x"2e098106",
   269 => x"8938810b",
   270 => x"fedc0c88",
   271 => x"c304800b",
   272 => x"fedc0c81",
   273 => x"5b807625",
   274 => x"80eb3878",
   275 => x"52765184",
   276 => x"812d80c1",
   277 => x"a452be88",
   278 => x"519ef02d",
   279 => x"bdec0880",
   280 => x"2ebc3880",
   281 => x"c1a45a83",
   282 => x"fc587970",
   283 => x"84055b08",
   284 => x"7083fe80",
   285 => x"0671882b",
   286 => x"83fe8006",
   287 => x"71882a07",
   288 => x"72882a83",
   289 => x"fe800673",
   290 => x"982a07fe",
   291 => x"c80cfec8",
   292 => x"0c56fc19",
   293 => x"59537780",
   294 => x"25d03889",
   295 => x"a504bdec",
   296 => x"085b8480",
   297 => x"56be8851",
   298 => x"9ec22dfc",
   299 => x"80168118",
   300 => x"585688c5",
   301 => x"047a5372",
   302 => x"bdec0c02",
   303 => x"ac050d04",
   304 => x"02fc050d",
   305 => x"ac962dfe",
   306 => x"c4518171",
   307 => x"0c82710c",
   308 => x"0284050d",
   309 => x"0402e805",
   310 => x"0d775680",
   311 => x"70565473",
   312 => x"7624b338",
   313 => x"80c7b408",
   314 => x"742eab38",
   315 => x"735199f8",
   316 => x"2dbdec08",
   317 => x"bdec0809",
   318 => x"810570bd",
   319 => x"ec08079f",
   320 => x"2a770581",
   321 => x"17575753",
   322 => x"53747624",
   323 => x"893880c7",
   324 => x"b4087426",
   325 => x"d73872bd",
   326 => x"ec0c0298",
   327 => x"050d0402",
   328 => x"fc050dbd",
   329 => x"98081351",
   330 => x"89d52dbd",
   331 => x"ec085187",
   332 => x"c22dbadc",
   333 => x"51adfa2d",
   334 => x"ac962d80",
   335 => x"5184e62d",
   336 => x"0284050d",
   337 => x"0402f405",
   338 => x"0d747678",
   339 => x"53545280",
   340 => x"71259738",
   341 => x"72708105",
   342 => x"5480f52d",
   343 => x"72708105",
   344 => x"5481b72d",
   345 => x"ff115170",
   346 => x"eb388072",
   347 => x"81b72d02",
   348 => x"8c050d04",
   349 => x"02dc050d",
   350 => x"80705a55",
   351 => x"74bd9808",
   352 => x"25b13880",
   353 => x"c7b40875",
   354 => x"2ea93878",
   355 => x"5199f82d",
   356 => x"bdec0809",
   357 => x"810570bd",
   358 => x"ec08079f",
   359 => x"2a760581",
   360 => x"1b5b5654",
   361 => x"74bd9808",
   362 => x"25893880",
   363 => x"c7b40879",
   364 => x"26d93880",
   365 => x"557880c7",
   366 => x"b4082781",
   367 => x"d0387851",
   368 => x"99f82dbd",
   369 => x"ec08802e",
   370 => x"81a538bd",
   371 => x"ec088b05",
   372 => x"80f52d70",
   373 => x"842a7081",
   374 => x"06771078",
   375 => x"842b80c5",
   376 => x"a40b80f5",
   377 => x"2d5c5c53",
   378 => x"51555673",
   379 => x"802e80c7",
   380 => x"38741682",
   381 => x"2b8db00b",
   382 => x"bbec120c",
   383 => x"54777531",
   384 => x"10be9c11",
   385 => x"55569074",
   386 => x"70810556",
   387 => x"81b72da0",
   388 => x"7481b72d",
   389 => x"7681ff06",
   390 => x"81165854",
   391 => x"73802e8a",
   392 => x"389c5380",
   393 => x"c5a4528c",
   394 => x"b0048b53",
   395 => x"bdec0852",
   396 => x"be9e1651",
   397 => x"8ce70474",
   398 => x"16822b8a",
   399 => x"9f0bbbec",
   400 => x"120c5476",
   401 => x"81ff0681",
   402 => x"16585473",
   403 => x"802e8a38",
   404 => x"9c5380c5",
   405 => x"a4528cdf",
   406 => x"048b53bd",
   407 => x"ec085277",
   408 => x"753110be",
   409 => x"9c055176",
   410 => x"558ac52d",
   411 => x"8d820474",
   412 => x"90297531",
   413 => x"7010be9c",
   414 => x"055154bd",
   415 => x"ec087481",
   416 => x"b72d8119",
   417 => x"59748b24",
   418 => x"a2388bb5",
   419 => x"04749029",
   420 => x"75317010",
   421 => x"be9c058c",
   422 => x"77315751",
   423 => x"54807481",
   424 => x"b72d9e14",
   425 => x"ff165654",
   426 => x"74f33802",
   427 => x"a4050d04",
   428 => x"02fc050d",
   429 => x"bd980813",
   430 => x"5189d52d",
   431 => x"bdec0880",
   432 => x"2e8838bd",
   433 => x"ec085192",
   434 => x"872d800b",
   435 => x"bd980c8a",
   436 => x"f42dacd9",
   437 => x"2d028405",
   438 => x"0d0402fc",
   439 => x"050d7251",
   440 => x"70fd2ead",
   441 => x"3870fd24",
   442 => x"8a3870fc",
   443 => x"2e80c438",
   444 => x"8ebb0470",
   445 => x"fe2eb138",
   446 => x"70ff2e09",
   447 => x"8106bc38",
   448 => x"bd980851",
   449 => x"70802eb3",
   450 => x"38ff11bd",
   451 => x"980c8ebb",
   452 => x"04bd9808",
   453 => x"f00570bd",
   454 => x"980c5170",
   455 => x"80259c38",
   456 => x"800bbd98",
   457 => x"0c8ebb04",
   458 => x"bd980881",
   459 => x"05bd980c",
   460 => x"8ebb04bd",
   461 => x"98089005",
   462 => x"bd980c8a",
   463 => x"f42dacd9",
   464 => x"2d028405",
   465 => x"0d0402fc",
   466 => x"050dbe94",
   467 => x"08fb06be",
   468 => x"940c7251",
   469 => x"8a9f2d02",
   470 => x"84050d04",
   471 => x"02fc050d",
   472 => x"be940884",
   473 => x"07be940c",
   474 => x"72518a9f",
   475 => x"2d028405",
   476 => x"0d0402fc",
   477 => x"050d800b",
   478 => x"bd980c8a",
   479 => x"f42dbbe4",
   480 => x"51adfa2d",
   481 => x"bbcc51ae",
   482 => x"8d2d0284",
   483 => x"050d0402",
   484 => x"f8050d80",
   485 => x"c8900882",
   486 => x"06bafc0b",
   487 => x"80f52d52",
   488 => x"5270802e",
   489 => x"85387181",
   490 => x"0752bb94",
   491 => x"0b80f52d",
   492 => x"5170802e",
   493 => x"85387184",
   494 => x"0752be98",
   495 => x"08802e85",
   496 => x"38719007",
   497 => x"5271bdec",
   498 => x"0c028805",
   499 => x"0d0402f4",
   500 => x"050d810b",
   501 => x"be980c90",
   502 => x"5186932d",
   503 => x"810bfec4",
   504 => x"0c900bfe",
   505 => x"c00c840b",
   506 => x"fec40c83",
   507 => x"0bfecc0c",
   508 => x"a9e22dab",
   509 => x"f72da9c5",
   510 => x"2da9c52d",
   511 => x"81f82d81",
   512 => x"5184e62d",
   513 => x"a9c52da9",
   514 => x"c52d8151",
   515 => x"84e62db8",
   516 => x"fc5185f2",
   517 => x"2d8452a3",
   518 => x"d02d939f",
   519 => x"2dbdec08",
   520 => x"802e8638",
   521 => x"fe5290b1",
   522 => x"04ff1252",
   523 => x"718024e7",
   524 => x"3871802e",
   525 => x"81833886",
   526 => x"c42db994",
   527 => x"5187c22d",
   528 => x"bdec0880",
   529 => x"2e8f38ba",
   530 => x"dc51adfa",
   531 => x"2d805184",
   532 => x"e62d90df",
   533 => x"04bdec08",
   534 => x"518ef22d",
   535 => x"ac832da9",
   536 => x"fb2dae93",
   537 => x"2dbdec08",
   538 => x"80c89408",
   539 => x"882b80c8",
   540 => x"980807fe",
   541 => x"d80c538f",
   542 => x"8f2dbdec",
   543 => x"08be9408",
   544 => x"2ea238bd",
   545 => x"ec08be94",
   546 => x"0cbdec08",
   547 => x"fec00c84",
   548 => x"52725184",
   549 => x"e62da9c5",
   550 => x"2da9c52d",
   551 => x"ff125271",
   552 => x"8025ee38",
   553 => x"72802e89",
   554 => x"388a0bfe",
   555 => x"c40c90df",
   556 => x"04820bfe",
   557 => x"c40c90df",
   558 => x"04b9a051",
   559 => x"85f22d80",
   560 => x"0bbdec0c",
   561 => x"028c050d",
   562 => x"0402e805",
   563 => x"0d77797b",
   564 => x"58555580",
   565 => x"53727625",
   566 => x"a3387470",
   567 => x"81055680",
   568 => x"f52d7470",
   569 => x"81055680",
   570 => x"f52d5252",
   571 => x"71712e86",
   572 => x"38815191",
   573 => x"fe048113",
   574 => x"5391d504",
   575 => x"805170bd",
   576 => x"ec0c0298",
   577 => x"050d0402",
   578 => x"ec050d76",
   579 => x"5574802e",
   580 => x"80da389a",
   581 => x"1580e02d",
   582 => x"51a88a2d",
   583 => x"bdec08bd",
   584 => x"ec0880c7",
   585 => x"d40cbdec",
   586 => x"08545480",
   587 => x"c7b00880",
   588 => x"2e993894",
   589 => x"1580e02d",
   590 => x"51a88a2d",
   591 => x"bdec0890",
   592 => x"2b83fff0",
   593 => x"0a067075",
   594 => x"07515372",
   595 => x"80c7d40c",
   596 => x"80c7a808",
   597 => x"fe147129",
   598 => x"80c7bc08",
   599 => x"0580c7d8",
   600 => x"0c70842b",
   601 => x"80c7b40c",
   602 => x"54939a04",
   603 => x"80c7c008",
   604 => x"80c7d40c",
   605 => x"80c7c408",
   606 => x"80c7d80c",
   607 => x"80c7b008",
   608 => x"802e8b38",
   609 => x"80c7a808",
   610 => x"842b5393",
   611 => x"950480c7",
   612 => x"c808842b",
   613 => x"537280c7",
   614 => x"b40c0294",
   615 => x"050d0402",
   616 => x"d8050d80",
   617 => x"0b80c7b0",
   618 => x"0c80c1a4",
   619 => x"528051a6",
   620 => x"ba2dbdec",
   621 => x"0854bdec",
   622 => x"088c38b9",
   623 => x"b45185f2",
   624 => x"2d735598",
   625 => x"fb048056",
   626 => x"810b80c7",
   627 => x"dc0c8853",
   628 => x"b9c05280",
   629 => x"c1da5191",
   630 => x"c92dbdec",
   631 => x"08762e09",
   632 => x"81068838",
   633 => x"bdec0880",
   634 => x"c7dc0c88",
   635 => x"53b9cc52",
   636 => x"80c1f651",
   637 => x"91c92dbd",
   638 => x"ec088838",
   639 => x"bdec0880",
   640 => x"c7dc0c80",
   641 => x"c7dc0880",
   642 => x"2e80fd38",
   643 => x"80c4ea0b",
   644 => x"80f52d80",
   645 => x"c4eb0b80",
   646 => x"f52d7198",
   647 => x"2b71902b",
   648 => x"0780c4ec",
   649 => x"0b80f52d",
   650 => x"70882b72",
   651 => x"0780c4ed",
   652 => x"0b80f52d",
   653 => x"710780c5",
   654 => x"a20b80f5",
   655 => x"2d80c5a3",
   656 => x"0b80f52d",
   657 => x"71882b07",
   658 => x"535f5452",
   659 => x"5a565755",
   660 => x"7381abaa",
   661 => x"2e098106",
   662 => x"8d387551",
   663 => x"a7da2dbd",
   664 => x"ec085694",
   665 => x"f3047382",
   666 => x"d4d52e87",
   667 => x"38b9d851",
   668 => x"95b80480",
   669 => x"c1a45275",
   670 => x"51a6ba2d",
   671 => x"bdec0855",
   672 => x"bdec0880",
   673 => x"2e83f438",
   674 => x"8853b9cc",
   675 => x"5280c1f6",
   676 => x"5191c92d",
   677 => x"bdec088a",
   678 => x"38810b80",
   679 => x"c7b00c95",
   680 => x"be048853",
   681 => x"b9c05280",
   682 => x"c1da5191",
   683 => x"c92dbdec",
   684 => x"08802e8a",
   685 => x"38b9ec51",
   686 => x"85f22d96",
   687 => x"9d0480c5",
   688 => x"a20b80f5",
   689 => x"2d547380",
   690 => x"d52e0981",
   691 => x"0680ce38",
   692 => x"80c5a30b",
   693 => x"80f52d54",
   694 => x"7381aa2e",
   695 => x"098106bd",
   696 => x"38800b80",
   697 => x"c1a40b80",
   698 => x"f52d5654",
   699 => x"7481e92e",
   700 => x"83388154",
   701 => x"7481eb2e",
   702 => x"8c388055",
   703 => x"73752e09",
   704 => x"810682f7",
   705 => x"3880c1af",
   706 => x"0b80f52d",
   707 => x"55748e38",
   708 => x"80c1b00b",
   709 => x"80f52d54",
   710 => x"73822e86",
   711 => x"38805598",
   712 => x"fb0480c1",
   713 => x"b10b80f5",
   714 => x"2d7080c7",
   715 => x"a80cff05",
   716 => x"80c7ac0c",
   717 => x"80c1b20b",
   718 => x"80f52d80",
   719 => x"c1b30b80",
   720 => x"f52d5876",
   721 => x"05778280",
   722 => x"29057080",
   723 => x"c7b80c80",
   724 => x"c1b40b80",
   725 => x"f52d7080",
   726 => x"c7cc0c80",
   727 => x"c7b00859",
   728 => x"57587680",
   729 => x"2e81b538",
   730 => x"8853b9cc",
   731 => x"5280c1f6",
   732 => x"5191c92d",
   733 => x"bdec0882",
   734 => x"823880c7",
   735 => x"a8087084",
   736 => x"2b80c7b4",
   737 => x"0c7080c7",
   738 => x"c80c80c1",
   739 => x"c90b80f5",
   740 => x"2d80c1c8",
   741 => x"0b80f52d",
   742 => x"71828029",
   743 => x"0580c1ca",
   744 => x"0b80f52d",
   745 => x"70848080",
   746 => x"291280c1",
   747 => x"cb0b80f5",
   748 => x"2d708180",
   749 => x"0a291270",
   750 => x"80c7d00c",
   751 => x"80c7cc08",
   752 => x"712980c7",
   753 => x"b8080570",
   754 => x"80c7bc0c",
   755 => x"80c1d10b",
   756 => x"80f52d80",
   757 => x"c1d00b80",
   758 => x"f52d7182",
   759 => x"80290580",
   760 => x"c1d20b80",
   761 => x"f52d7084",
   762 => x"80802912",
   763 => x"80c1d30b",
   764 => x"80f52d70",
   765 => x"982b81f0",
   766 => x"0a067205",
   767 => x"7080c7c0",
   768 => x"0cfe117e",
   769 => x"29770580",
   770 => x"c7c40c52",
   771 => x"59524354",
   772 => x"5e515259",
   773 => x"525d5759",
   774 => x"5798f404",
   775 => x"80c1b60b",
   776 => x"80f52d80",
   777 => x"c1b50b80",
   778 => x"f52d7182",
   779 => x"80290570",
   780 => x"80c7b40c",
   781 => x"70a02983",
   782 => x"ff057089",
   783 => x"2a7080c7",
   784 => x"c80c80c1",
   785 => x"bb0b80f5",
   786 => x"2d80c1ba",
   787 => x"0b80f52d",
   788 => x"71828029",
   789 => x"057080c7",
   790 => x"d00c7b71",
   791 => x"291e7080",
   792 => x"c7c40c7d",
   793 => x"80c7c00c",
   794 => x"730580c7",
   795 => x"bc0c555e",
   796 => x"51515555",
   797 => x"80519287",
   798 => x"2d815574",
   799 => x"bdec0c02",
   800 => x"a8050d04",
   801 => x"02ec050d",
   802 => x"7670872c",
   803 => x"7180ff06",
   804 => x"55565480",
   805 => x"c7b0088a",
   806 => x"3873882c",
   807 => x"7481ff06",
   808 => x"545580c1",
   809 => x"a45280c7",
   810 => x"b8081551",
   811 => x"a6ba2dbd",
   812 => x"ec0854bd",
   813 => x"ec08802e",
   814 => x"b63880c7",
   815 => x"b008802e",
   816 => x"99387284",
   817 => x"2980c1a4",
   818 => x"05700852",
   819 => x"53a7da2d",
   820 => x"bdec08f0",
   821 => x"0a065399",
   822 => x"ed047210",
   823 => x"80c1a405",
   824 => x"7080e02d",
   825 => x"5253a88a",
   826 => x"2dbdec08",
   827 => x"53725473",
   828 => x"bdec0c02",
   829 => x"94050d04",
   830 => x"02e0050d",
   831 => x"7970842c",
   832 => x"80c7d808",
   833 => x"05718f06",
   834 => x"52555372",
   835 => x"8a3880c1",
   836 => x"a4527351",
   837 => x"a6ba2d72",
   838 => x"a02980c1",
   839 => x"a4055480",
   840 => x"7480f52d",
   841 => x"56537473",
   842 => x"2e833881",
   843 => x"537481e5",
   844 => x"2e81f138",
   845 => x"81707406",
   846 => x"54587280",
   847 => x"2e81e538",
   848 => x"8b1480f5",
   849 => x"2d70832a",
   850 => x"79065856",
   851 => x"769938bd",
   852 => x"9c085372",
   853 => x"89387280",
   854 => x"c5a40b81",
   855 => x"b72d76bd",
   856 => x"9c0c7353",
   857 => x"9ca60475",
   858 => x"8f2e0981",
   859 => x"0681b538",
   860 => x"749f068d",
   861 => x"2980c597",
   862 => x"11515381",
   863 => x"1480f52d",
   864 => x"73708105",
   865 => x"5581b72d",
   866 => x"831480f5",
   867 => x"2d737081",
   868 => x"055581b7",
   869 => x"2d851480",
   870 => x"f52d7370",
   871 => x"81055581",
   872 => x"b72d8714",
   873 => x"80f52d73",
   874 => x"70810555",
   875 => x"81b72d89",
   876 => x"1480f52d",
   877 => x"73708105",
   878 => x"5581b72d",
   879 => x"8e1480f5",
   880 => x"2d737081",
   881 => x"055581b7",
   882 => x"2d901480",
   883 => x"f52d7370",
   884 => x"81055581",
   885 => x"b72d9214",
   886 => x"80f52d73",
   887 => x"70810555",
   888 => x"81b72d94",
   889 => x"1480f52d",
   890 => x"73708105",
   891 => x"5581b72d",
   892 => x"961480f5",
   893 => x"2d737081",
   894 => x"055581b7",
   895 => x"2d981480",
   896 => x"f52d7370",
   897 => x"81055581",
   898 => x"b72d9c14",
   899 => x"80f52d73",
   900 => x"70810555",
   901 => x"81b72d9e",
   902 => x"1480f52d",
   903 => x"7381b72d",
   904 => x"77bd9c0c",
   905 => x"805372bd",
   906 => x"ec0c02a0",
   907 => x"050d0402",
   908 => x"cc050d7e",
   909 => x"605e5a80",
   910 => x"0b80c7d4",
   911 => x"0880c7d8",
   912 => x"08595c56",
   913 => x"805880c7",
   914 => x"b408782e",
   915 => x"81b23877",
   916 => x"8f06a017",
   917 => x"57547391",
   918 => x"3880c1a4",
   919 => x"52765181",
   920 => x"1757a6ba",
   921 => x"2d80c1a4",
   922 => x"56807680",
   923 => x"f52d5654",
   924 => x"74742e83",
   925 => x"38815474",
   926 => x"81e52e80",
   927 => x"f7388170",
   928 => x"7506555c",
   929 => x"73802e80",
   930 => x"eb388b16",
   931 => x"80f52d98",
   932 => x"06597880",
   933 => x"df388b53",
   934 => x"7c527551",
   935 => x"91c92dbd",
   936 => x"ec0880d0",
   937 => x"389c1608",
   938 => x"51a7da2d",
   939 => x"bdec0884",
   940 => x"1b0c9a16",
   941 => x"80e02d51",
   942 => x"a88a2dbd",
   943 => x"ec08bdec",
   944 => x"08881c0c",
   945 => x"bdec0855",
   946 => x"5580c7b0",
   947 => x"08802e98",
   948 => x"38941680",
   949 => x"e02d51a8",
   950 => x"8a2dbdec",
   951 => x"08902b83",
   952 => x"fff00a06",
   953 => x"70165154",
   954 => x"73881b0c",
   955 => x"787a0c7b",
   956 => x"549eb904",
   957 => x"81185880",
   958 => x"c7b40878",
   959 => x"26fed038",
   960 => x"80c7b008",
   961 => x"802eb038",
   962 => x"7a519984",
   963 => x"2dbdec08",
   964 => x"bdec0880",
   965 => x"fffffff8",
   966 => x"06555b73",
   967 => x"80ffffff",
   968 => x"f82e9438",
   969 => x"bdec08fe",
   970 => x"0580c7a8",
   971 => x"082980c7",
   972 => x"bc080557",
   973 => x"9cc40480",
   974 => x"5473bdec",
   975 => x"0c02b405",
   976 => x"0d0402f4",
   977 => x"050d7470",
   978 => x"08810571",
   979 => x"0c700880",
   980 => x"c7ac0806",
   981 => x"5353718e",
   982 => x"38881308",
   983 => x"5199842d",
   984 => x"bdec0888",
   985 => x"140c810b",
   986 => x"bdec0c02",
   987 => x"8c050d04",
   988 => x"02f0050d",
   989 => x"75881108",
   990 => x"fe0580c7",
   991 => x"a8082980",
   992 => x"c7bc0811",
   993 => x"720880c7",
   994 => x"ac080605",
   995 => x"79555354",
   996 => x"54a6ba2d",
   997 => x"0290050d",
   998 => x"0402f005",
   999 => x"0d758811",
  1000 => x"08fe0580",
  1001 => x"c7a80829",
  1002 => x"80c7bc08",
  1003 => x"11720880",
  1004 => x"c7ac0806",
  1005 => x"05795553",
  1006 => x"5454a4fa",
  1007 => x"2d029005",
  1008 => x"0d0402f4",
  1009 => x"050dd452",
  1010 => x"81ff720c",
  1011 => x"71085381",
  1012 => x"ff720c72",
  1013 => x"882b83fe",
  1014 => x"80067208",
  1015 => x"7081ff06",
  1016 => x"51525381",
  1017 => x"ff720c72",
  1018 => x"7107882b",
  1019 => x"72087081",
  1020 => x"ff065152",
  1021 => x"5381ff72",
  1022 => x"0c727107",
  1023 => x"882b7208",
  1024 => x"7081ff06",
  1025 => x"7207bdec",
  1026 => x"0c525302",
  1027 => x"8c050d04",
  1028 => x"02f4050d",
  1029 => x"74767181",
  1030 => x"ff06d40c",
  1031 => x"535380c7",
  1032 => x"e0088538",
  1033 => x"71892b52",
  1034 => x"71982ad4",
  1035 => x"0c71902a",
  1036 => x"7081ff06",
  1037 => x"d40c5171",
  1038 => x"882a7081",
  1039 => x"ff06d40c",
  1040 => x"517181ff",
  1041 => x"06d40c72",
  1042 => x"902a7081",
  1043 => x"ff06d40c",
  1044 => x"51d40870",
  1045 => x"81ff0651",
  1046 => x"5182b8bf",
  1047 => x"527081ff",
  1048 => x"2e098106",
  1049 => x"943881ff",
  1050 => x"0bd40cd4",
  1051 => x"087081ff",
  1052 => x"06ff1454",
  1053 => x"515171e5",
  1054 => x"3870bdec",
  1055 => x"0c028c05",
  1056 => x"0d0402fc",
  1057 => x"050d81c7",
  1058 => x"5181ff0b",
  1059 => x"d40cff11",
  1060 => x"51708025",
  1061 => x"f4380284",
  1062 => x"050d0402",
  1063 => x"f0050da1",
  1064 => x"822d8fcf",
  1065 => x"53805287",
  1066 => x"fc80f751",
  1067 => x"a0902dbd",
  1068 => x"ec0854bd",
  1069 => x"ec08812e",
  1070 => x"098106a3",
  1071 => x"3881ff0b",
  1072 => x"d40c820a",
  1073 => x"52849c80",
  1074 => x"e951a090",
  1075 => x"2dbdec08",
  1076 => x"8b3881ff",
  1077 => x"0bd40c73",
  1078 => x"53a1e504",
  1079 => x"a1822dff",
  1080 => x"135372c1",
  1081 => x"3872bdec",
  1082 => x"0c029005",
  1083 => x"0d0402f4",
  1084 => x"050d81ff",
  1085 => x"0bd40c93",
  1086 => x"53805287",
  1087 => x"fc80c151",
  1088 => x"a0902dbd",
  1089 => x"ec088b38",
  1090 => x"81ff0bd4",
  1091 => x"0c8153a2",
  1092 => x"9b04a182",
  1093 => x"2dff1353",
  1094 => x"72df3872",
  1095 => x"bdec0c02",
  1096 => x"8c050d04",
  1097 => x"02f0050d",
  1098 => x"a1822d83",
  1099 => x"aa52849c",
  1100 => x"80c851a0",
  1101 => x"902dbdec",
  1102 => x"08812e09",
  1103 => x"81069238",
  1104 => x"9fc22dbd",
  1105 => x"ec0883ff",
  1106 => x"ff065372",
  1107 => x"83aa2e97",
  1108 => x"38a1ee2d",
  1109 => x"a2e20481",
  1110 => x"54a3c704",
  1111 => x"b9f85185",
  1112 => x"f22d8054",
  1113 => x"a3c70481",
  1114 => x"ff0bd40c",
  1115 => x"b153a19b",
  1116 => x"2dbdec08",
  1117 => x"802e80c0",
  1118 => x"38805287",
  1119 => x"fc80fa51",
  1120 => x"a0902dbd",
  1121 => x"ec08b138",
  1122 => x"81ff0bd4",
  1123 => x"0cd40853",
  1124 => x"81ff0bd4",
  1125 => x"0c81ff0b",
  1126 => x"d40c81ff",
  1127 => x"0bd40c81",
  1128 => x"ff0bd40c",
  1129 => x"72862a70",
  1130 => x"8106bdec",
  1131 => x"08565153",
  1132 => x"72802e93",
  1133 => x"38a2d704",
  1134 => x"72822eff",
  1135 => x"9f38ff13",
  1136 => x"5372ffaa",
  1137 => x"38725473",
  1138 => x"bdec0c02",
  1139 => x"90050d04",
  1140 => x"02f0050d",
  1141 => x"810b80c7",
  1142 => x"e00c8454",
  1143 => x"d008708f",
  1144 => x"2a708106",
  1145 => x"51515372",
  1146 => x"f33872d0",
  1147 => x"0ca1822d",
  1148 => x"ba885185",
  1149 => x"f22dd008",
  1150 => x"708f2a70",
  1151 => x"81065151",
  1152 => x"5372f338",
  1153 => x"810bd00c",
  1154 => x"b1538052",
  1155 => x"84d480c0",
  1156 => x"51a0902d",
  1157 => x"bdec0881",
  1158 => x"2ea13872",
  1159 => x"822e0981",
  1160 => x"068c38ba",
  1161 => x"945185f2",
  1162 => x"2d8053a4",
  1163 => x"f104ff13",
  1164 => x"5372d738",
  1165 => x"ff145473",
  1166 => x"ffa238a2",
  1167 => x"a42dbdec",
  1168 => x"0880c7e0",
  1169 => x"0cbdec08",
  1170 => x"8b388152",
  1171 => x"87fc80d0",
  1172 => x"51a0902d",
  1173 => x"81ff0bd4",
  1174 => x"0cd00870",
  1175 => x"8f2a7081",
  1176 => x"06515153",
  1177 => x"72f33872",
  1178 => x"d00c81ff",
  1179 => x"0bd40c81",
  1180 => x"5372bdec",
  1181 => x"0c029005",
  1182 => x"0d0402e8",
  1183 => x"050d7856",
  1184 => x"81ff0bd4",
  1185 => x"0cd00870",
  1186 => x"8f2a7081",
  1187 => x"06515153",
  1188 => x"72f33882",
  1189 => x"810bd00c",
  1190 => x"81ff0bd4",
  1191 => x"0c775287",
  1192 => x"fc80d851",
  1193 => x"a0902dbd",
  1194 => x"ec08802e",
  1195 => x"8c38baac",
  1196 => x"5185f22d",
  1197 => x"8153a6b1",
  1198 => x"0481ff0b",
  1199 => x"d40c81fe",
  1200 => x"0bd40c80",
  1201 => x"ff557570",
  1202 => x"84055708",
  1203 => x"70982ad4",
  1204 => x"0c70902c",
  1205 => x"7081ff06",
  1206 => x"d40c5470",
  1207 => x"882c7081",
  1208 => x"ff06d40c",
  1209 => x"547081ff",
  1210 => x"06d40c54",
  1211 => x"ff155574",
  1212 => x"8025d338",
  1213 => x"81ff0bd4",
  1214 => x"0c81ff0b",
  1215 => x"d40c81ff",
  1216 => x"0bd40c86",
  1217 => x"8da05481",
  1218 => x"ff0bd40c",
  1219 => x"d40881ff",
  1220 => x"06557487",
  1221 => x"38ff1454",
  1222 => x"73ed3881",
  1223 => x"ff0bd40c",
  1224 => x"d008708f",
  1225 => x"2a708106",
  1226 => x"51515372",
  1227 => x"f33872d0",
  1228 => x"0c72bdec",
  1229 => x"0c029805",
  1230 => x"0d0402e8",
  1231 => x"050d7855",
  1232 => x"805681ff",
  1233 => x"0bd40cd0",
  1234 => x"08708f2a",
  1235 => x"70810651",
  1236 => x"515372f3",
  1237 => x"3882810b",
  1238 => x"d00c81ff",
  1239 => x"0bd40c77",
  1240 => x"5287fc80",
  1241 => x"d151a090",
  1242 => x"2d80dbc6",
  1243 => x"df54bdec",
  1244 => x"08802e8a",
  1245 => x"38babc51",
  1246 => x"85f22da7",
  1247 => x"d10481ff",
  1248 => x"0bd40cd4",
  1249 => x"087081ff",
  1250 => x"06515372",
  1251 => x"81fe2e09",
  1252 => x"81069d38",
  1253 => x"80ff539f",
  1254 => x"c22dbdec",
  1255 => x"08757084",
  1256 => x"05570cff",
  1257 => x"13537280",
  1258 => x"25ed3881",
  1259 => x"56a7b604",
  1260 => x"ff145473",
  1261 => x"c93881ff",
  1262 => x"0bd40c81",
  1263 => x"ff0bd40c",
  1264 => x"d008708f",
  1265 => x"2a708106",
  1266 => x"51515372",
  1267 => x"f33872d0",
  1268 => x"0c75bdec",
  1269 => x"0c029805",
  1270 => x"0d0402f4",
  1271 => x"050d7470",
  1272 => x"882a83fe",
  1273 => x"80067072",
  1274 => x"982a0772",
  1275 => x"882b87fc",
  1276 => x"80800673",
  1277 => x"982b81f0",
  1278 => x"0a067173",
  1279 => x"0707bdec",
  1280 => x"0c565153",
  1281 => x"51028c05",
  1282 => x"0d0402f8",
  1283 => x"050d028e",
  1284 => x"0580f52d",
  1285 => x"74882b07",
  1286 => x"7083ffff",
  1287 => x"06bdec0c",
  1288 => x"51028805",
  1289 => x"0d0402fc",
  1290 => x"050d7251",
  1291 => x"80710c80",
  1292 => x"0b84120c",
  1293 => x"0284050d",
  1294 => x"0402f005",
  1295 => x"0d757008",
  1296 => x"84120853",
  1297 => x"5353ff54",
  1298 => x"71712ea8",
  1299 => x"38abfd2d",
  1300 => x"84130870",
  1301 => x"84291488",
  1302 => x"11700870",
  1303 => x"81ff0684",
  1304 => x"18088111",
  1305 => x"8706841a",
  1306 => x"0c535155",
  1307 => x"515151ab",
  1308 => x"f72d7154",
  1309 => x"73bdec0c",
  1310 => x"0290050d",
  1311 => x"0402f805",
  1312 => x"0dabfd2d",
  1313 => x"e008708b",
  1314 => x"2a708106",
  1315 => x"51525270",
  1316 => x"802ea138",
  1317 => x"80c7e408",
  1318 => x"70842980",
  1319 => x"c7ec0573",
  1320 => x"81ff0671",
  1321 => x"0c515180",
  1322 => x"c7e40881",
  1323 => x"11870680",
  1324 => x"c7e40c51",
  1325 => x"800b80c8",
  1326 => x"8c0cabf0",
  1327 => x"2dabf72d",
  1328 => x"0288050d",
  1329 => x"0402fc05",
  1330 => x"0dabfd2d",
  1331 => x"810b80c8",
  1332 => x"8c0cabf7",
  1333 => x"2d80c88c",
  1334 => x"085170f9",
  1335 => x"38028405",
  1336 => x"0d0402fc",
  1337 => x"050d80c7",
  1338 => x"e451a8a6",
  1339 => x"2da8fd51",
  1340 => x"abec2dab",
  1341 => x"962d0284",
  1342 => x"050d0402",
  1343 => x"f4050daa",
  1344 => x"fd04bdec",
  1345 => x"0881f02e",
  1346 => x"09810689",
  1347 => x"38810bbd",
  1348 => x"e00caafd",
  1349 => x"04bdec08",
  1350 => x"81e02e09",
  1351 => x"81068938",
  1352 => x"810bbde4",
  1353 => x"0caafd04",
  1354 => x"bdec0852",
  1355 => x"bde40880",
  1356 => x"2e8838bd",
  1357 => x"ec088180",
  1358 => x"05527184",
  1359 => x"2c728f06",
  1360 => x"5353bde0",
  1361 => x"08802e99",
  1362 => x"38728429",
  1363 => x"bda00572",
  1364 => x"1381712b",
  1365 => x"70097308",
  1366 => x"06730c51",
  1367 => x"5353aaf3",
  1368 => x"04728429",
  1369 => x"bda00572",
  1370 => x"1383712b",
  1371 => x"72080772",
  1372 => x"0c535380",
  1373 => x"0bbde40c",
  1374 => x"800bbde0",
  1375 => x"0c80c7e4",
  1376 => x"51a8b92d",
  1377 => x"bdec08ff",
  1378 => x"24fef738",
  1379 => x"800bbdec",
  1380 => x"0c028c05",
  1381 => x"0d0402f8",
  1382 => x"050dbda0",
  1383 => x"528f5180",
  1384 => x"72708405",
  1385 => x"540cff11",
  1386 => x"51708025",
  1387 => x"f2380288",
  1388 => x"050d0402",
  1389 => x"f0050d75",
  1390 => x"51abfd2d",
  1391 => x"70822cfc",
  1392 => x"06bda011",
  1393 => x"72109e06",
  1394 => x"71087072",
  1395 => x"2a708306",
  1396 => x"82742b70",
  1397 => x"09740676",
  1398 => x"0c545156",
  1399 => x"57535153",
  1400 => x"abf72d71",
  1401 => x"bdec0c02",
  1402 => x"90050d04",
  1403 => x"71980c04",
  1404 => x"ffb008bd",
  1405 => x"ec0c0481",
  1406 => x"0bffb00c",
  1407 => x"04800bff",
  1408 => x"b00c0402",
  1409 => x"fc050d81",
  1410 => x"0bbde80c",
  1411 => x"815184e6",
  1412 => x"2d028405",
  1413 => x"0d0402fc",
  1414 => x"050d800b",
  1415 => x"bde80c80",
  1416 => x"5184e62d",
  1417 => x"0284050d",
  1418 => x"0402ec05",
  1419 => x"0d765480",
  1420 => x"52870b88",
  1421 => x"1580f52d",
  1422 => x"56537472",
  1423 => x"248338a0",
  1424 => x"53725182",
  1425 => x"ef2d8112",
  1426 => x"8b1580f5",
  1427 => x"2d545272",
  1428 => x"7225de38",
  1429 => x"0294050d",
  1430 => x"0402f005",
  1431 => x"0d80c89c",
  1432 => x"085481f8",
  1433 => x"2d800b80",
  1434 => x"c8a00c73",
  1435 => x"08802e81",
  1436 => x"8438820b",
  1437 => x"be800c80",
  1438 => x"c8a0088f",
  1439 => x"06bdfc0c",
  1440 => x"73085271",
  1441 => x"832e9638",
  1442 => x"71832689",
  1443 => x"3871812e",
  1444 => x"af38adde",
  1445 => x"0471852e",
  1446 => x"9f38adde",
  1447 => x"04881480",
  1448 => x"f52d8415",
  1449 => x"08bacc53",
  1450 => x"545285f2",
  1451 => x"2d718429",
  1452 => x"13700852",
  1453 => x"52ade204",
  1454 => x"7351aca9",
  1455 => x"2dadde04",
  1456 => x"80c89008",
  1457 => x"8815082c",
  1458 => x"70810651",
  1459 => x"5271802e",
  1460 => x"8738bad0",
  1461 => x"51addb04",
  1462 => x"bad45185",
  1463 => x"f22d8414",
  1464 => x"085185f2",
  1465 => x"2d80c8a0",
  1466 => x"08810580",
  1467 => x"c8a00c8c",
  1468 => x"1454aceb",
  1469 => x"04029005",
  1470 => x"0d047180",
  1471 => x"c89c0cac",
  1472 => x"d92d80c8",
  1473 => x"a008ff05",
  1474 => x"80c8a40c",
  1475 => x"047180c8",
  1476 => x"a80c0402",
  1477 => x"e8050d80",
  1478 => x"c89c0880",
  1479 => x"c8a80857",
  1480 => x"5580f851",
  1481 => x"abb32dbd",
  1482 => x"ec08812a",
  1483 => x"70810651",
  1484 => x"52719b38",
  1485 => x"8751abb3",
  1486 => x"2dbdec08",
  1487 => x"812a7081",
  1488 => x"06515271",
  1489 => x"802eb138",
  1490 => x"aece04a9",
  1491 => x"fb2d8751",
  1492 => x"abb32dbd",
  1493 => x"ec08f438",
  1494 => x"aede04a9",
  1495 => x"fb2d80f8",
  1496 => x"51abb32d",
  1497 => x"bdec08f3",
  1498 => x"38bde808",
  1499 => x"813270bd",
  1500 => x"e80c7052",
  1501 => x"5284e62d",
  1502 => x"800b80c8",
  1503 => x"940c800b",
  1504 => x"80c8980c",
  1505 => x"bde80882",
  1506 => x"fd3880da",
  1507 => x"51abb32d",
  1508 => x"bdec0880",
  1509 => x"2e8c3880",
  1510 => x"c8940881",
  1511 => x"800780c8",
  1512 => x"940c80d9",
  1513 => x"51abb32d",
  1514 => x"bdec0880",
  1515 => x"2e8c3880",
  1516 => x"c8940880",
  1517 => x"c00780c8",
  1518 => x"940c8194",
  1519 => x"51abb32d",
  1520 => x"bdec0880",
  1521 => x"2e8b3880",
  1522 => x"c8940890",
  1523 => x"0780c894",
  1524 => x"0c819151",
  1525 => x"abb32dbd",
  1526 => x"ec08802e",
  1527 => x"8b3880c8",
  1528 => x"9408a007",
  1529 => x"80c8940c",
  1530 => x"81f551ab",
  1531 => x"b32dbdec",
  1532 => x"08802e8b",
  1533 => x"3880c894",
  1534 => x"08810780",
  1535 => x"c8940c81",
  1536 => x"f251abb3",
  1537 => x"2dbdec08",
  1538 => x"802e8b38",
  1539 => x"80c89408",
  1540 => x"820780c8",
  1541 => x"940c81eb",
  1542 => x"51abb32d",
  1543 => x"bdec0880",
  1544 => x"2e8b3880",
  1545 => x"c8940884",
  1546 => x"0780c894",
  1547 => x"0c81f451",
  1548 => x"abb32dbd",
  1549 => x"ec08802e",
  1550 => x"8b3880c8",
  1551 => x"94088807",
  1552 => x"80c8940c",
  1553 => x"80d851ab",
  1554 => x"b32dbdec",
  1555 => x"08802e8c",
  1556 => x"3880c898",
  1557 => x"08818007",
  1558 => x"80c8980c",
  1559 => x"9251abb3",
  1560 => x"2dbdec08",
  1561 => x"802e8c38",
  1562 => x"80c89808",
  1563 => x"80c00780",
  1564 => x"c8980c94",
  1565 => x"51abb32d",
  1566 => x"bdec0880",
  1567 => x"2e8b3880",
  1568 => x"c8980890",
  1569 => x"0780c898",
  1570 => x"0c9151ab",
  1571 => x"b32dbdec",
  1572 => x"08802e8b",
  1573 => x"3880c898",
  1574 => x"08a00780",
  1575 => x"c8980c9d",
  1576 => x"51abb32d",
  1577 => x"bdec0880",
  1578 => x"2e8b3880",
  1579 => x"c8980881",
  1580 => x"0780c898",
  1581 => x"0c9b51ab",
  1582 => x"b32dbdec",
  1583 => x"08802e8b",
  1584 => x"3880c898",
  1585 => x"08820780",
  1586 => x"c8980c9c",
  1587 => x"51abb32d",
  1588 => x"bdec0880",
  1589 => x"2e8b3880",
  1590 => x"c8980884",
  1591 => x"0780c898",
  1592 => x"0ca351ab",
  1593 => x"b32dbdec",
  1594 => x"08802e8b",
  1595 => x"3880c898",
  1596 => x"08880780",
  1597 => x"c8980c81",
  1598 => x"fd51abb3",
  1599 => x"2d81fa51",
  1600 => x"abb32db7",
  1601 => x"ce0481f5",
  1602 => x"51abb32d",
  1603 => x"bdec0881",
  1604 => x"2a708106",
  1605 => x"51527180",
  1606 => x"2eb33880",
  1607 => x"c8a40852",
  1608 => x"71802e8a",
  1609 => x"38ff1280",
  1610 => x"c8a40cb2",
  1611 => x"cd0480c8",
  1612 => x"a0081080",
  1613 => x"c8a00805",
  1614 => x"70842916",
  1615 => x"51528812",
  1616 => x"08802e89",
  1617 => x"38ff5188",
  1618 => x"12085271",
  1619 => x"2d81f251",
  1620 => x"abb32dbd",
  1621 => x"ec08812a",
  1622 => x"70810651",
  1623 => x"5271802e",
  1624 => x"b43880c8",
  1625 => x"a008ff11",
  1626 => x"80c8a408",
  1627 => x"56535373",
  1628 => x"72258a38",
  1629 => x"811480c8",
  1630 => x"a40cb395",
  1631 => x"04721013",
  1632 => x"70842916",
  1633 => x"51528812",
  1634 => x"08802e89",
  1635 => x"38fe5188",
  1636 => x"12085271",
  1637 => x"2d81fd51",
  1638 => x"abb32dbd",
  1639 => x"ec08812a",
  1640 => x"70810651",
  1641 => x"5271802e",
  1642 => x"b13880c8",
  1643 => x"a408802e",
  1644 => x"8a38800b",
  1645 => x"80c8a40c",
  1646 => x"b3da0480",
  1647 => x"c8a00810",
  1648 => x"80c8a008",
  1649 => x"05708429",
  1650 => x"16515288",
  1651 => x"1208802e",
  1652 => x"8938fd51",
  1653 => x"88120852",
  1654 => x"712d81fa",
  1655 => x"51abb32d",
  1656 => x"bdec0881",
  1657 => x"2a708106",
  1658 => x"51527180",
  1659 => x"2eb13880",
  1660 => x"c8a008ff",
  1661 => x"11545280",
  1662 => x"c8a40873",
  1663 => x"25893872",
  1664 => x"80c8a40c",
  1665 => x"b49f0471",
  1666 => x"10127084",
  1667 => x"29165152",
  1668 => x"88120880",
  1669 => x"2e8938fc",
  1670 => x"51881208",
  1671 => x"52712d80",
  1672 => x"c8a40870",
  1673 => x"53547380",
  1674 => x"2e8a388c",
  1675 => x"15ff1555",
  1676 => x"55b4a604",
  1677 => x"820bbe80",
  1678 => x"0c718f06",
  1679 => x"bdfc0c81",
  1680 => x"eb51abb3",
  1681 => x"2dbdec08",
  1682 => x"812a7081",
  1683 => x"06515271",
  1684 => x"802ead38",
  1685 => x"7408852e",
  1686 => x"098106a4",
  1687 => x"38881580",
  1688 => x"f52dff05",
  1689 => x"52718816",
  1690 => x"81b72d71",
  1691 => x"982b5271",
  1692 => x"80258838",
  1693 => x"800b8816",
  1694 => x"81b72d74",
  1695 => x"51aca92d",
  1696 => x"81f451ab",
  1697 => x"b32dbdec",
  1698 => x"08812a70",
  1699 => x"81065152",
  1700 => x"71802eb3",
  1701 => x"38740885",
  1702 => x"2e098106",
  1703 => x"aa388815",
  1704 => x"80f52d81",
  1705 => x"05527188",
  1706 => x"1681b72d",
  1707 => x"7181ff06",
  1708 => x"8b1680f5",
  1709 => x"2d545272",
  1710 => x"72278738",
  1711 => x"72881681",
  1712 => x"b72d7451",
  1713 => x"aca92d80",
  1714 => x"da51abb3",
  1715 => x"2dbdec08",
  1716 => x"812a7081",
  1717 => x"06515271",
  1718 => x"802e81ac",
  1719 => x"3880c89c",
  1720 => x"0880c8a4",
  1721 => x"08555373",
  1722 => x"802e8a38",
  1723 => x"8c13ff15",
  1724 => x"5553b5e7",
  1725 => x"04720852",
  1726 => x"71822ea6",
  1727 => x"38718226",
  1728 => x"89387181",
  1729 => x"2eaa38b7",
  1730 => x"88047183",
  1731 => x"2eb43871",
  1732 => x"842e0981",
  1733 => x"0680f138",
  1734 => x"88130851",
  1735 => x"adfa2db7",
  1736 => x"880480c8",
  1737 => x"a4085188",
  1738 => x"13085271",
  1739 => x"2db78804",
  1740 => x"810b8814",
  1741 => x"082b80c8",
  1742 => x"90083280",
  1743 => x"c8900cb6",
  1744 => x"dd048813",
  1745 => x"80f52d81",
  1746 => x"058b1480",
  1747 => x"f52d5354",
  1748 => x"71742483",
  1749 => x"38805473",
  1750 => x"881481b7",
  1751 => x"2dacd92d",
  1752 => x"b7880475",
  1753 => x"08802ea3",
  1754 => x"38750851",
  1755 => x"abb32dbd",
  1756 => x"ec088106",
  1757 => x"5271802e",
  1758 => x"8c3880c8",
  1759 => x"a4085184",
  1760 => x"16085271",
  1761 => x"2d881656",
  1762 => x"75d93880",
  1763 => x"54800bbe",
  1764 => x"800c738f",
  1765 => x"06bdfc0c",
  1766 => x"a0527380",
  1767 => x"c8a4082e",
  1768 => x"09810699",
  1769 => x"3880c8a0",
  1770 => x"08ff0574",
  1771 => x"32700981",
  1772 => x"05707207",
  1773 => x"9f2a9171",
  1774 => x"31515153",
  1775 => x"53715182",
  1776 => x"ef2d8114",
  1777 => x"548e7425",
  1778 => x"c438bde8",
  1779 => x"085271bd",
  1780 => x"ec0c0298",
  1781 => x"050d0400",
  1782 => x"00ffffff",
  1783 => x"ff00ffff",
  1784 => x"ffff00ff",
  1785 => x"ffffff00",
  1786 => x"52657365",
  1787 => x"74000000",
  1788 => x"53617665",
  1789 => x"20736574",
  1790 => x"74696e67",
  1791 => x"73000000",
  1792 => x"5363616e",
  1793 => x"6c696e65",
  1794 => x"73000000",
  1795 => x"4c6f6164",
  1796 => x"20524f4d",
  1797 => x"20100000",
  1798 => x"45786974",
  1799 => x"00000000",
  1800 => x"50432045",
  1801 => x"6e67696e",
  1802 => x"65206d6f",
  1803 => x"64650000",
  1804 => x"54757262",
  1805 => x"6f677261",
  1806 => x"66782031",
  1807 => x"36206d6f",
  1808 => x"64650000",
  1809 => x"56474120",
  1810 => x"2d203331",
  1811 => x"4b487a2c",
  1812 => x"20363048",
  1813 => x"7a000000",
  1814 => x"5456202d",
  1815 => x"20343830",
  1816 => x"692c2036",
  1817 => x"30487a00",
  1818 => x"4261636b",
  1819 => x"00000000",
  1820 => x"46504741",
  1821 => x"50434520",
  1822 => x"43464700",
  1823 => x"496e6974",
  1824 => x"69616c69",
  1825 => x"7a696e67",
  1826 => x"20534420",
  1827 => x"63617264",
  1828 => x"0a000000",
  1829 => x"424f4f54",
  1830 => x"20202020",
  1831 => x"50434500",
  1832 => x"43617264",
  1833 => x"20696e69",
  1834 => x"74206661",
  1835 => x"696c6564",
  1836 => x"0a000000",
  1837 => x"4d425220",
  1838 => x"6661696c",
  1839 => x"0a000000",
  1840 => x"46415431",
  1841 => x"36202020",
  1842 => x"00000000",
  1843 => x"46415433",
  1844 => x"32202020",
  1845 => x"00000000",
  1846 => x"4e6f2070",
  1847 => x"61727469",
  1848 => x"74696f6e",
  1849 => x"20736967",
  1850 => x"0a000000",
  1851 => x"42616420",
  1852 => x"70617274",
  1853 => x"0a000000",
  1854 => x"53444843",
  1855 => x"20657272",
  1856 => x"6f72210a",
  1857 => x"00000000",
  1858 => x"53442069",
  1859 => x"6e69742e",
  1860 => x"2e2e0a00",
  1861 => x"53442063",
  1862 => x"61726420",
  1863 => x"72657365",
  1864 => x"74206661",
  1865 => x"696c6564",
  1866 => x"210a0000",
  1867 => x"57726974",
  1868 => x"65206661",
  1869 => x"696c6564",
  1870 => x"0a000000",
  1871 => x"52656164",
  1872 => x"20666169",
  1873 => x"6c65640a",
  1874 => x"00000000",
  1875 => x"16200000",
  1876 => x"14200000",
  1877 => x"15200000",
  1878 => x"00000002",
  1879 => x"00000002",
  1880 => x"00001be8",
  1881 => x"000004c0",
  1882 => x"00000002",
  1883 => x"00001bf0",
  1884 => x"0000037d",
  1885 => x"00000003",
  1886 => x"00001dc4",
  1887 => x"00000002",
  1888 => x"00000001",
  1889 => x"00001c00",
  1890 => x"00000001",
  1891 => x"00000003",
  1892 => x"00001dbc",
  1893 => x"00000002",
  1894 => x"00000002",
  1895 => x"00001c0c",
  1896 => x"00000772",
  1897 => x"00000002",
  1898 => x"00001c18",
  1899 => x"00001616",
  1900 => x"00000000",
  1901 => x"00000000",
  1902 => x"00000000",
  1903 => x"00001c20",
  1904 => x"00001c30",
  1905 => x"00001c44",
  1906 => x"00001c58",
  1907 => x"0000004d",
  1908 => x"00000746",
  1909 => x"0000002c",
  1910 => x"0000075c",
  1911 => x"00000000",
  1912 => x"00000000",
  1913 => x"00000002",
  1914 => x"00001f1c",
  1915 => x"0000051f",
  1916 => x"00000002",
  1917 => x"00001f3a",
  1918 => x"0000051f",
  1919 => x"00000002",
  1920 => x"00001f58",
  1921 => x"0000051f",
  1922 => x"00000002",
  1923 => x"00001f76",
  1924 => x"0000051f",
  1925 => x"00000002",
  1926 => x"00001f94",
  1927 => x"0000051f",
  1928 => x"00000002",
  1929 => x"00001fb2",
  1930 => x"0000051f",
  1931 => x"00000002",
  1932 => x"00001fd0",
  1933 => x"0000051f",
  1934 => x"00000002",
  1935 => x"00001fee",
  1936 => x"0000051f",
  1937 => x"00000002",
  1938 => x"0000200c",
  1939 => x"0000051f",
  1940 => x"00000002",
  1941 => x"0000202a",
  1942 => x"0000051f",
  1943 => x"00000002",
  1944 => x"00002048",
  1945 => x"0000051f",
  1946 => x"00000002",
  1947 => x"00002066",
  1948 => x"0000051f",
  1949 => x"00000002",
  1950 => x"00002084",
  1951 => x"0000051f",
  1952 => x"00000004",
  1953 => x"00001c68",
  1954 => x"00001d5c",
  1955 => x"00000000",
  1956 => x"00000000",
  1957 => x"000006da",
  1958 => x"00000000",
  1959 => x"00000000",
  1960 => x"00000000",
  1961 => x"00000000",
  1962 => x"00000000",
  1963 => x"00000000",
  1964 => x"00000000",
  1965 => x"00000000",
  1966 => x"00000000",
  1967 => x"00000000",
  1968 => x"00000000",
  1969 => x"00000000",
  1970 => x"00000000",
  1971 => x"00000000",
  1972 => x"00000000",
  1973 => x"00000000",
  1974 => x"00000000",
  1975 => x"00000000",
  1976 => x"00000000",
  1977 => x"00000000",
  1978 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

