-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb6",
     9 => x"b4080b0b",
    10 => x"0bb6b808",
    11 => x"0b0b0bb6",
    12 => x"bc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b6bc0c0b",
    16 => x"0b0bb6b8",
    17 => x"0c0b0b0b",
    18 => x"b6b40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb0a4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b6b470bd",
    57 => x"b0278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8d8c0402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b6c40c9f",
    65 => x"0bb6c80c",
    66 => x"a0717081",
    67 => x"055334b6",
    68 => x"c808ff05",
    69 => x"b6c80cb6",
    70 => x"c8088025",
    71 => x"eb38b6c4",
    72 => x"08ff05b6",
    73 => x"c40cb6c4",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb6c4",
    94 => x"08258f38",
    95 => x"82b22db6",
    96 => x"c408ff05",
    97 => x"b6c40c82",
    98 => x"f404b6c4",
    99 => x"08b6c808",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b6c408",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b6",
   108 => x"c8088105",
   109 => x"b6c80cb6",
   110 => x"c808519f",
   111 => x"7125e238",
   112 => x"800bb6c8",
   113 => x"0cb6c408",
   114 => x"8105b6c4",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b6c80881",
   120 => x"05b6c80c",
   121 => x"b6c808a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b6c80cb6",
   125 => x"c4088105",
   126 => x"b6c40c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb6",
   155 => x"cc0cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb6cc",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b6cc0884",
   167 => x"07b6cc0c",
   168 => x"5573842b",
   169 => x"87e87125",
   170 => x"83713170",
   171 => x"0b0b0bb3",
   172 => x"a40c8171",
   173 => x"2bf6880c",
   174 => x"fea413ff",
   175 => x"122c7888",
   176 => x"29ff9405",
   177 => x"70812cb6",
   178 => x"cc085258",
   179 => x"52555152",
   180 => x"5476802e",
   181 => x"85387081",
   182 => x"075170f6",
   183 => x"940c7109",
   184 => x"8105f680",
   185 => x"0c720981",
   186 => x"05f6840c",
   187 => x"0294050d",
   188 => x"0402f405",
   189 => x"0d745372",
   190 => x"70810554",
   191 => x"80f52d52",
   192 => x"71802e89",
   193 => x"38715182",
   194 => x"ee2d85f7",
   195 => x"04028c05",
   196 => x"0d0402f4",
   197 => x"050d7470",
   198 => x"8206bd94",
   199 => x"0cb3c071",
   200 => x"81065454",
   201 => x"51718814",
   202 => x"81b72d70",
   203 => x"822a7081",
   204 => x"06515170",
   205 => x"a01481b7",
   206 => x"2d70b6b4",
   207 => x"0c028c05",
   208 => x"0d0402f8",
   209 => x"050db1bc",
   210 => x"52b6d051",
   211 => x"96aa2db6",
   212 => x"b408802e",
   213 => x"9d38b8b4",
   214 => x"52b6d051",
   215 => x"98e02db8",
   216 => x"b408b6dc",
   217 => x"0cb8b408",
   218 => x"fec00cb8",
   219 => x"b4085186",
   220 => x"922d0288",
   221 => x"050d0402",
   222 => x"f0050db1",
   223 => x"bc52b6d0",
   224 => x"5196aa2d",
   225 => x"b6b40880",
   226 => x"2ea538b6",
   227 => x"dc08b8b4",
   228 => x"0cb8b854",
   229 => x"80fd5380",
   230 => x"74708405",
   231 => x"560cff13",
   232 => x"53728025",
   233 => x"f238b8b4",
   234 => x"52b6d051",
   235 => x"99862d02",
   236 => x"90050d04",
   237 => x"02d4050d",
   238 => x"b6dc08fe",
   239 => x"c00c810b",
   240 => x"fec40c84",
   241 => x"0bfec40c",
   242 => x"7c52b6d0",
   243 => x"5196aa2d",
   244 => x"b6b40853",
   245 => x"b6b40880",
   246 => x"2e81cc38",
   247 => x"b6d40856",
   248 => x"800bff17",
   249 => x"58597679",
   250 => x"2e8b3881",
   251 => x"1977812a",
   252 => x"585976f7",
   253 => x"38f71976",
   254 => x"9fff0654",
   255 => x"5972802e",
   256 => x"8b38fc80",
   257 => x"16b6d052",
   258 => x"5698b32d",
   259 => x"75b08080",
   260 => x"2e098106",
   261 => x"8938820b",
   262 => x"fedc0c88",
   263 => x"b5047598",
   264 => x"80802e09",
   265 => x"81068938",
   266 => x"810bfedc",
   267 => x"0c88b504",
   268 => x"800bfedc",
   269 => x"0c815b80",
   270 => x"762580e9",
   271 => x"38785276",
   272 => x"5184802d",
   273 => x"b8b452b6",
   274 => x"d05198e0",
   275 => x"2db6b408",
   276 => x"802ebb38",
   277 => x"b8b45a83",
   278 => x"fc587970",
   279 => x"84055b08",
   280 => x"7083fe80",
   281 => x"0671882b",
   282 => x"83fe8006",
   283 => x"71882a07",
   284 => x"72882a83",
   285 => x"fe800673",
   286 => x"982a07fe",
   287 => x"c80cfec8",
   288 => x"0c56fc19",
   289 => x"59537780",
   290 => x"25d03889",
   291 => x"9504b6b4",
   292 => x"085b8480",
   293 => x"56b6d051",
   294 => x"98b32dfc",
   295 => x"80168118",
   296 => x"585688b7",
   297 => x"047a5372",
   298 => x"b6b40c02",
   299 => x"ac050d04",
   300 => x"02fc050d",
   301 => x"a5f42dfe",
   302 => x"c4518171",
   303 => x"0c82710c",
   304 => x"0284050d",
   305 => x"0402f405",
   306 => x"0d741015",
   307 => x"708429b4",
   308 => x"b4057008",
   309 => x"55515272",
   310 => x"802e9038",
   311 => x"7280f52d",
   312 => x"5271802e",
   313 => x"86387251",
   314 => x"87b42db3",
   315 => x"a851a7d2",
   316 => x"2da5f42d",
   317 => x"805184e5",
   318 => x"2d028c05",
   319 => x"0d0402e8",
   320 => x"050d8070",
   321 => x"565675b5",
   322 => x"e40825af",
   323 => x"38bcc008",
   324 => x"762ea838",
   325 => x"745195d5",
   326 => x"2db6b408",
   327 => x"09810570",
   328 => x"b6b40807",
   329 => x"9f2a7705",
   330 => x"81175757",
   331 => x"5275b5e4",
   332 => x"08258838",
   333 => x"bcc00875",
   334 => x"26da3880",
   335 => x"5674bcc0",
   336 => x"082780d0",
   337 => x"38745195",
   338 => x"d52d7584",
   339 => x"2b52b6b4",
   340 => x"08802eae",
   341 => x"38b6e412",
   342 => x"8117b6b4",
   343 => x"08565752",
   344 => x"8a537370",
   345 => x"81055580",
   346 => x"f52d7270",
   347 => x"81055481",
   348 => x"b72dff13",
   349 => x"53728025",
   350 => x"e9388072",
   351 => x"81b72d8b",
   352 => x"8b04b6b4",
   353 => x"08b6e413",
   354 => x"81b72d81",
   355 => x"15558b76",
   356 => x"25ffaa38",
   357 => x"0298050d",
   358 => x"0402fc05",
   359 => x"0d725170",
   360 => x"fd2ead38",
   361 => x"70fd248a",
   362 => x"3870fc2e",
   363 => x"80c4388b",
   364 => x"fa0470fe",
   365 => x"2eb13870",
   366 => x"ff2e0981",
   367 => x"06bc38b5",
   368 => x"e4085170",
   369 => x"802eb338",
   370 => x"ff11b5e4",
   371 => x"0c8bfa04",
   372 => x"b5e408f0",
   373 => x"0570b5e4",
   374 => x"0c517080",
   375 => x"259c3880",
   376 => x"0bb5e40c",
   377 => x"8bfa04b5",
   378 => x"e4088105",
   379 => x"b5e40c8b",
   380 => x"fa04b5e4",
   381 => x"089005b5",
   382 => x"e40c89fe",
   383 => x"2da6b72d",
   384 => x"0284050d",
   385 => x"0402fc05",
   386 => x"0db6dc08",
   387 => x"fb06b6dc",
   388 => x"0c725189",
   389 => x"c52d0284",
   390 => x"050d0402",
   391 => x"fc050db6",
   392 => x"dc088407",
   393 => x"b6dc0c72",
   394 => x"5189c52d",
   395 => x"0284050d",
   396 => x"0402fc05",
   397 => x"0d800bb5",
   398 => x"e40c89fe",
   399 => x"2db4b051",
   400 => x"a7d22db4",
   401 => x"9851a7e2",
   402 => x"2d028405",
   403 => x"0d0402f8",
   404 => x"050dbd94",
   405 => x"088206b3",
   406 => x"c80b80f5",
   407 => x"2d525270",
   408 => x"802e8538",
   409 => x"71810752",
   410 => x"b3e00b80",
   411 => x"f52d5170",
   412 => x"802e8538",
   413 => x"71840752",
   414 => x"b6e00880",
   415 => x"2e853871",
   416 => x"90075271",
   417 => x"b6b40c02",
   418 => x"88050d04",
   419 => x"02f4050d",
   420 => x"810bb6e0",
   421 => x"0c905186",
   422 => x"922d810b",
   423 => x"fec40c90",
   424 => x"0bfec00c",
   425 => x"840bfec4",
   426 => x"0c830bfe",
   427 => x"cc0ca3c2",
   428 => x"2da5d52d",
   429 => x"a3a72da3",
   430 => x"a72d81f7",
   431 => x"2d815184",
   432 => x"e52da3a7",
   433 => x"2da3a72d",
   434 => x"815184e5",
   435 => x"2db1c851",
   436 => x"85f12d84",
   437 => x"529db92d",
   438 => x"8fc32db6",
   439 => x"b408802e",
   440 => x"8638fe52",
   441 => x"8def04ff",
   442 => x"12527180",
   443 => x"24e73871",
   444 => x"802e8181",
   445 => x"3886c22d",
   446 => x"b1e05187",
   447 => x"b42db6b4",
   448 => x"08802e8f",
   449 => x"38b3a851",
   450 => x"a7d22d80",
   451 => x"5184e52d",
   452 => x"8e9d04b6",
   453 => x"b408518c",
   454 => x"b12da5e1",
   455 => x"2da3da2d",
   456 => x"a7e72db6",
   457 => x"b408bd98",
   458 => x"08882bbd",
   459 => x"9c0807fe",
   460 => x"d80c538c",
   461 => x"ce2db6b4",
   462 => x"08b6dc08",
   463 => x"2ea238b6",
   464 => x"b408b6dc",
   465 => x"0cb6b408",
   466 => x"fec00c84",
   467 => x"52725184",
   468 => x"e52da3a7",
   469 => x"2da3a72d",
   470 => x"ff125271",
   471 => x"8025ee38",
   472 => x"72802e89",
   473 => x"388a0bfe",
   474 => x"c40c8e9d",
   475 => x"04820bfe",
   476 => x"c40c8e9d",
   477 => x"04b1ec51",
   478 => x"85f12d80",
   479 => x"0bb6b40c",
   480 => x"028c050d",
   481 => x"0402e805",
   482 => x"0d77797b",
   483 => x"58555580",
   484 => x"53727625",
   485 => x"a3387470",
   486 => x"81055680",
   487 => x"f52d7470",
   488 => x"81055680",
   489 => x"f52d5252",
   490 => x"71712e86",
   491 => x"3881518f",
   492 => x"ba048113",
   493 => x"538f9104",
   494 => x"805170b6",
   495 => x"b40c0298",
   496 => x"050d0402",
   497 => x"d8050d80",
   498 => x"0bbcbc0c",
   499 => x"b8b45280",
   500 => x"51a0a12d",
   501 => x"b6b40854",
   502 => x"b6b4088c",
   503 => x"38b28051",
   504 => x"85f12d73",
   505 => x"5594de04",
   506 => x"8056810b",
   507 => x"bce00c88",
   508 => x"53b28c52",
   509 => x"b8ea518f",
   510 => x"852db6b4",
   511 => x"08762e09",
   512 => x"81068738",
   513 => x"b6b408bc",
   514 => x"e00c8853",
   515 => x"b29852b9",
   516 => x"86518f85",
   517 => x"2db6b408",
   518 => x"8738b6b4",
   519 => x"08bce00c",
   520 => x"bce00880",
   521 => x"2e80f638",
   522 => x"bbfa0b80",
   523 => x"f52dbbfb",
   524 => x"0b80f52d",
   525 => x"71982b71",
   526 => x"902b07bb",
   527 => x"fc0b80f5",
   528 => x"2d70882b",
   529 => x"7207bbfd",
   530 => x"0b80f52d",
   531 => x"7107bcb2",
   532 => x"0b80f52d",
   533 => x"bcb30b80",
   534 => x"f52d7188",
   535 => x"2b07535f",
   536 => x"54525a56",
   537 => x"57557381",
   538 => x"abaa2e09",
   539 => x"81068d38",
   540 => x"7551a1c1",
   541 => x"2db6b408",
   542 => x"56918904",
   543 => x"7382d4d5",
   544 => x"2e8738b2",
   545 => x"a45191ca",
   546 => x"04b8b452",
   547 => x"7551a0a1",
   548 => x"2db6b408",
   549 => x"55b6b408",
   550 => x"802e83c2",
   551 => x"388853b2",
   552 => x"9852b986",
   553 => x"518f852d",
   554 => x"b6b40889",
   555 => x"38810bbc",
   556 => x"bc0c91d0",
   557 => x"048853b2",
   558 => x"8c52b8ea",
   559 => x"518f852d",
   560 => x"b6b40880",
   561 => x"2e8a38b2",
   562 => x"b85185f1",
   563 => x"2d92aa04",
   564 => x"bcb20b80",
   565 => x"f52d5473",
   566 => x"80d52e09",
   567 => x"810680ca",
   568 => x"38bcb30b",
   569 => x"80f52d54",
   570 => x"7381aa2e",
   571 => x"098106ba",
   572 => x"38800bb8",
   573 => x"b40b80f5",
   574 => x"2d565474",
   575 => x"81e92e83",
   576 => x"38815474",
   577 => x"81eb2e8c",
   578 => x"38805573",
   579 => x"752e0981",
   580 => x"0682cb38",
   581 => x"b8bf0b80",
   582 => x"f52d5574",
   583 => x"8d38b8c0",
   584 => x"0b80f52d",
   585 => x"5473822e",
   586 => x"86388055",
   587 => x"94de04b8",
   588 => x"c10b80f5",
   589 => x"2d70bcb4",
   590 => x"0cff05bc",
   591 => x"b80cb8c2",
   592 => x"0b80f52d",
   593 => x"b8c30b80",
   594 => x"f52d5876",
   595 => x"05778280",
   596 => x"290570bc",
   597 => x"c40cb8c4",
   598 => x"0b80f52d",
   599 => x"70bcd80c",
   600 => x"bcbc0859",
   601 => x"57587680",
   602 => x"2e81a338",
   603 => x"8853b298",
   604 => x"52b98651",
   605 => x"8f852db6",
   606 => x"b40881e2",
   607 => x"38bcb408",
   608 => x"70842bbc",
   609 => x"c00c70bc",
   610 => x"d40cb8d9",
   611 => x"0b80f52d",
   612 => x"b8d80b80",
   613 => x"f52d7182",
   614 => x"802905b8",
   615 => x"da0b80f5",
   616 => x"2d708480",
   617 => x"802912b8",
   618 => x"db0b80f5",
   619 => x"2d708180",
   620 => x"0a291270",
   621 => x"bcdc0cbc",
   622 => x"d8087129",
   623 => x"bcc40805",
   624 => x"70bcc80c",
   625 => x"b8e10b80",
   626 => x"f52db8e0",
   627 => x"0b80f52d",
   628 => x"71828029",
   629 => x"05b8e20b",
   630 => x"80f52d70",
   631 => x"84808029",
   632 => x"12b8e30b",
   633 => x"80f52d70",
   634 => x"982b81f0",
   635 => x"0a067205",
   636 => x"70bccc0c",
   637 => x"fe117e29",
   638 => x"7705bcd0",
   639 => x"0c525952",
   640 => x"43545e51",
   641 => x"5259525d",
   642 => x"57595794",
   643 => x"dc04b8c6",
   644 => x"0b80f52d",
   645 => x"b8c50b80",
   646 => x"f52d7182",
   647 => x"80290570",
   648 => x"bcc00c70",
   649 => x"a02983ff",
   650 => x"0570892a",
   651 => x"70bcd40c",
   652 => x"b8cb0b80",
   653 => x"f52db8ca",
   654 => x"0b80f52d",
   655 => x"71828029",
   656 => x"0570bcdc",
   657 => x"0c7b7129",
   658 => x"1e70bcd0",
   659 => x"0c7dbccc",
   660 => x"0c7305bc",
   661 => x"c80c555e",
   662 => x"51515555",
   663 => x"815574b6",
   664 => x"b40c02a8",
   665 => x"050d0402",
   666 => x"ec050d76",
   667 => x"70872c71",
   668 => x"80ff0655",
   669 => x"5654bcbc",
   670 => x"088a3873",
   671 => x"882c7481",
   672 => x"ff065455",
   673 => x"b8b452bc",
   674 => x"c4081551",
   675 => x"a0a12db6",
   676 => x"b40854b6",
   677 => x"b408802e",
   678 => x"b338bcbc",
   679 => x"08802e98",
   680 => x"38728429",
   681 => x"b8b40570",
   682 => x"085253a1",
   683 => x"c12db6b4",
   684 => x"08f00a06",
   685 => x"5395ca04",
   686 => x"7210b8b4",
   687 => x"057080e0",
   688 => x"2d5253a1",
   689 => x"f12db6b4",
   690 => x"08537254",
   691 => x"73b6b40c",
   692 => x"0294050d",
   693 => x"0402ec05",
   694 => x"0d767084",
   695 => x"2cbcd008",
   696 => x"05718f06",
   697 => x"52555372",
   698 => x"8938b8b4",
   699 => x"527351a0",
   700 => x"a12d72a0",
   701 => x"29b8b405",
   702 => x"54807480",
   703 => x"f52d5455",
   704 => x"72752e83",
   705 => x"38815572",
   706 => x"81e52e93",
   707 => x"3874802e",
   708 => x"8e388b14",
   709 => x"80f52d98",
   710 => x"06537280",
   711 => x"2e833880",
   712 => x"5473b6b4",
   713 => x"0c029405",
   714 => x"0d0402cc",
   715 => x"050d7e60",
   716 => x"5e5a800b",
   717 => x"bccc08bc",
   718 => x"d008595c",
   719 => x"568058bc",
   720 => x"c008782e",
   721 => x"81ae3877",
   722 => x"8f06a017",
   723 => x"5754738f",
   724 => x"38b8b452",
   725 => x"76518117",
   726 => x"57a0a12d",
   727 => x"b8b45680",
   728 => x"7680f52d",
   729 => x"56547474",
   730 => x"2e833881",
   731 => x"547481e5",
   732 => x"2e80f638",
   733 => x"81707506",
   734 => x"555c7380",
   735 => x"2e80ea38",
   736 => x"8b1680f5",
   737 => x"2d980659",
   738 => x"7880de38",
   739 => x"8b537c52",
   740 => x"75518f85",
   741 => x"2db6b408",
   742 => x"80cf389c",
   743 => x"160851a1",
   744 => x"c12db6b4",
   745 => x"08841b0c",
   746 => x"9a1680e0",
   747 => x"2d51a1f1",
   748 => x"2db6b408",
   749 => x"b6b40888",
   750 => x"1c0cb6b4",
   751 => x"085555bc",
   752 => x"bc08802e",
   753 => x"98389416",
   754 => x"80e02d51",
   755 => x"a1f12db6",
   756 => x"b408902b",
   757 => x"83fff00a",
   758 => x"06701651",
   759 => x"5473881b",
   760 => x"0c787a0c",
   761 => x"7b5498aa",
   762 => x"04811858",
   763 => x"bcc00878",
   764 => x"26fed438",
   765 => x"bcbc0880",
   766 => x"2eae387a",
   767 => x"5194e72d",
   768 => x"b6b408b6",
   769 => x"b40880ff",
   770 => x"fffff806",
   771 => x"555b7380",
   772 => x"fffffff8",
   773 => x"2e9238b6",
   774 => x"b408fe05",
   775 => x"bcb40829",
   776 => x"bcc80805",
   777 => x"5796bd04",
   778 => x"805473b6",
   779 => x"b40c02b4",
   780 => x"050d0402",
   781 => x"f4050d74",
   782 => x"70088105",
   783 => x"710c7008",
   784 => x"bcb80806",
   785 => x"5353718e",
   786 => x"38881308",
   787 => x"5194e72d",
   788 => x"b6b40888",
   789 => x"140c810b",
   790 => x"b6b40c02",
   791 => x"8c050d04",
   792 => x"02f0050d",
   793 => x"75881108",
   794 => x"fe05bcb4",
   795 => x"0829bcc8",
   796 => x"08117208",
   797 => x"bcb80806",
   798 => x"05795553",
   799 => x"5454a0a1",
   800 => x"2d029005",
   801 => x"0d0402f0",
   802 => x"050d7588",
   803 => x"1108fe05",
   804 => x"bcb40829",
   805 => x"bcc80811",
   806 => x"7208bcb8",
   807 => x"08060579",
   808 => x"55535454",
   809 => x"9ee12d02",
   810 => x"90050d04",
   811 => x"02f4050d",
   812 => x"d45281ff",
   813 => x"720c7108",
   814 => x"5381ff72",
   815 => x"0c72882b",
   816 => x"83fe8006",
   817 => x"72087081",
   818 => x"ff065152",
   819 => x"5381ff72",
   820 => x"0c727107",
   821 => x"882b7208",
   822 => x"7081ff06",
   823 => x"51525381",
   824 => x"ff720c72",
   825 => x"7107882b",
   826 => x"72087081",
   827 => x"ff067207",
   828 => x"b6b40c52",
   829 => x"53028c05",
   830 => x"0d0402f4",
   831 => x"050d7476",
   832 => x"7181ff06",
   833 => x"d40c5353",
   834 => x"bce40885",
   835 => x"3871892b",
   836 => x"5271982a",
   837 => x"d40c7190",
   838 => x"2a7081ff",
   839 => x"06d40c51",
   840 => x"71882a70",
   841 => x"81ff06d4",
   842 => x"0c517181",
   843 => x"ff06d40c",
   844 => x"72902a70",
   845 => x"81ff06d4",
   846 => x"0c51d408",
   847 => x"7081ff06",
   848 => x"515182b8",
   849 => x"bf527081",
   850 => x"ff2e0981",
   851 => x"06943881",
   852 => x"ff0bd40c",
   853 => x"d4087081",
   854 => x"ff06ff14",
   855 => x"54515171",
   856 => x"e53870b6",
   857 => x"b40c028c",
   858 => x"050d0402",
   859 => x"fc050d81",
   860 => x"c75181ff",
   861 => x"0bd40cff",
   862 => x"11517080",
   863 => x"25f43802",
   864 => x"84050d04",
   865 => x"02f0050d",
   866 => x"9aeb2d8f",
   867 => x"cf538052",
   868 => x"87fc80f7",
   869 => x"5199fa2d",
   870 => x"b6b40854",
   871 => x"b6b40881",
   872 => x"2e098106",
   873 => x"a33881ff",
   874 => x"0bd40c82",
   875 => x"0a52849c",
   876 => x"80e95199",
   877 => x"fa2db6b4",
   878 => x"088b3881",
   879 => x"ff0bd40c",
   880 => x"73539bce",
   881 => x"049aeb2d",
   882 => x"ff135372",
   883 => x"c13872b6",
   884 => x"b40c0290",
   885 => x"050d0402",
   886 => x"f4050d81",
   887 => x"ff0bd40c",
   888 => x"93538052",
   889 => x"87fc80c1",
   890 => x"5199fa2d",
   891 => x"b6b4088b",
   892 => x"3881ff0b",
   893 => x"d40c8153",
   894 => x"9c84049a",
   895 => x"eb2dff13",
   896 => x"5372df38",
   897 => x"72b6b40c",
   898 => x"028c050d",
   899 => x"0402f005",
   900 => x"0d9aeb2d",
   901 => x"83aa5284",
   902 => x"9c80c851",
   903 => x"99fa2db6",
   904 => x"b408812e",
   905 => x"09810692",
   906 => x"3899ac2d",
   907 => x"b6b40883",
   908 => x"ffff0653",
   909 => x"7283aa2e",
   910 => x"97389bd7",
   911 => x"2d9ccb04",
   912 => x"81549db0",
   913 => x"04b2c451",
   914 => x"85f12d80",
   915 => x"549db004",
   916 => x"81ff0bd4",
   917 => x"0cb1539b",
   918 => x"842db6b4",
   919 => x"08802e80",
   920 => x"c0388052",
   921 => x"87fc80fa",
   922 => x"5199fa2d",
   923 => x"b6b408b1",
   924 => x"3881ff0b",
   925 => x"d40cd408",
   926 => x"5381ff0b",
   927 => x"d40c81ff",
   928 => x"0bd40c81",
   929 => x"ff0bd40c",
   930 => x"81ff0bd4",
   931 => x"0c72862a",
   932 => x"708106b6",
   933 => x"b4085651",
   934 => x"5372802e",
   935 => x"93389cc0",
   936 => x"0472822e",
   937 => x"ff9f38ff",
   938 => x"135372ff",
   939 => x"aa387254",
   940 => x"73b6b40c",
   941 => x"0290050d",
   942 => x"0402f005",
   943 => x"0d810bbc",
   944 => x"e40c8454",
   945 => x"d008708f",
   946 => x"2a708106",
   947 => x"51515372",
   948 => x"f33872d0",
   949 => x"0c9aeb2d",
   950 => x"b2d45185",
   951 => x"f12dd008",
   952 => x"708f2a70",
   953 => x"81065151",
   954 => x"5372f338",
   955 => x"810bd00c",
   956 => x"b1538052",
   957 => x"84d480c0",
   958 => x"5199fa2d",
   959 => x"b6b40881",
   960 => x"2ea13872",
   961 => x"822e0981",
   962 => x"068c38b2",
   963 => x"e05185f1",
   964 => x"2d80539e",
   965 => x"d804ff13",
   966 => x"5372d738",
   967 => x"ff145473",
   968 => x"ffa2389c",
   969 => x"8d2db6b4",
   970 => x"08bce40c",
   971 => x"b6b4088b",
   972 => x"38815287",
   973 => x"fc80d051",
   974 => x"99fa2d81",
   975 => x"ff0bd40c",
   976 => x"d008708f",
   977 => x"2a708106",
   978 => x"51515372",
   979 => x"f33872d0",
   980 => x"0c81ff0b",
   981 => x"d40c8153",
   982 => x"72b6b40c",
   983 => x"0290050d",
   984 => x"0402e805",
   985 => x"0d785681",
   986 => x"ff0bd40c",
   987 => x"d008708f",
   988 => x"2a708106",
   989 => x"51515372",
   990 => x"f3388281",
   991 => x"0bd00c81",
   992 => x"ff0bd40c",
   993 => x"775287fc",
   994 => x"80d85199",
   995 => x"fa2db6b4",
   996 => x"08802e8c",
   997 => x"38b2f851",
   998 => x"85f12d81",
   999 => x"53a09804",
  1000 => x"81ff0bd4",
  1001 => x"0c81fe0b",
  1002 => x"d40c80ff",
  1003 => x"55757084",
  1004 => x"05570870",
  1005 => x"982ad40c",
  1006 => x"70902c70",
  1007 => x"81ff06d4",
  1008 => x"0c547088",
  1009 => x"2c7081ff",
  1010 => x"06d40c54",
  1011 => x"7081ff06",
  1012 => x"d40c54ff",
  1013 => x"15557480",
  1014 => x"25d33881",
  1015 => x"ff0bd40c",
  1016 => x"81ff0bd4",
  1017 => x"0c81ff0b",
  1018 => x"d40c868d",
  1019 => x"a05481ff",
  1020 => x"0bd40cd4",
  1021 => x"0881ff06",
  1022 => x"55748738",
  1023 => x"ff145473",
  1024 => x"ed3881ff",
  1025 => x"0bd40cd0",
  1026 => x"08708f2a",
  1027 => x"70810651",
  1028 => x"515372f3",
  1029 => x"3872d00c",
  1030 => x"72b6b40c",
  1031 => x"0298050d",
  1032 => x"0402e805",
  1033 => x"0d785580",
  1034 => x"5681ff0b",
  1035 => x"d40cd008",
  1036 => x"708f2a70",
  1037 => x"81065151",
  1038 => x"5372f338",
  1039 => x"82810bd0",
  1040 => x"0c81ff0b",
  1041 => x"d40c7752",
  1042 => x"87fc80d1",
  1043 => x"5199fa2d",
  1044 => x"80dbc6df",
  1045 => x"54b6b408",
  1046 => x"802e8a38",
  1047 => x"b3885185",
  1048 => x"f12da1b8",
  1049 => x"0481ff0b",
  1050 => x"d40cd408",
  1051 => x"7081ff06",
  1052 => x"51537281",
  1053 => x"fe2e0981",
  1054 => x"069d3880",
  1055 => x"ff5399ac",
  1056 => x"2db6b408",
  1057 => x"75708405",
  1058 => x"570cff13",
  1059 => x"53728025",
  1060 => x"ed388156",
  1061 => x"a19d04ff",
  1062 => x"145473c9",
  1063 => x"3881ff0b",
  1064 => x"d40c81ff",
  1065 => x"0bd40cd0",
  1066 => x"08708f2a",
  1067 => x"70810651",
  1068 => x"515372f3",
  1069 => x"3872d00c",
  1070 => x"75b6b40c",
  1071 => x"0298050d",
  1072 => x"0402f405",
  1073 => x"0d747088",
  1074 => x"2a83fe80",
  1075 => x"06707298",
  1076 => x"2a077288",
  1077 => x"2b87fc80",
  1078 => x"80067398",
  1079 => x"2b81f00a",
  1080 => x"06717307",
  1081 => x"07b6b40c",
  1082 => x"56515351",
  1083 => x"028c050d",
  1084 => x"0402f805",
  1085 => x"0d028e05",
  1086 => x"80f52d74",
  1087 => x"882b0770",
  1088 => x"83ffff06",
  1089 => x"b6b40c51",
  1090 => x"0288050d",
  1091 => x"0402fc05",
  1092 => x"0d725180",
  1093 => x"710c800b",
  1094 => x"84120c02",
  1095 => x"84050d04",
  1096 => x"02f0050d",
  1097 => x"75700884",
  1098 => x"12085353",
  1099 => x"53ff5471",
  1100 => x"712ea838",
  1101 => x"a5db2d84",
  1102 => x"13087084",
  1103 => x"29148811",
  1104 => x"70087081",
  1105 => x"ff068418",
  1106 => x"08811187",
  1107 => x"06841a0c",
  1108 => x"53515551",
  1109 => x"5151a5d5",
  1110 => x"2d715473",
  1111 => x"b6b40c02",
  1112 => x"90050d04",
  1113 => x"02f8050d",
  1114 => x"a5db2de0",
  1115 => x"08708b2a",
  1116 => x"70810651",
  1117 => x"52527080",
  1118 => x"2e9d38bc",
  1119 => x"e8087084",
  1120 => x"29bcf005",
  1121 => x"7381ff06",
  1122 => x"710c5151",
  1123 => x"bce80881",
  1124 => x"118706bc",
  1125 => x"e80c5180",
  1126 => x"0bbd900c",
  1127 => x"a5ce2da5",
  1128 => x"d52d0288",
  1129 => x"050d0402",
  1130 => x"fc050da5",
  1131 => x"db2d810b",
  1132 => x"bd900ca5",
  1133 => x"d52dbd90",
  1134 => x"085170fa",
  1135 => x"38028405",
  1136 => x"0d0402fc",
  1137 => x"050dbce8",
  1138 => x"51a28d2d",
  1139 => x"a2e451a5",
  1140 => x"ca2da4f4",
  1141 => x"2d028405",
  1142 => x"0d0402f4",
  1143 => x"050da4dc",
  1144 => x"04b6b408",
  1145 => x"81f02e09",
  1146 => x"81068938",
  1147 => x"810bb6a8",
  1148 => x"0ca4dc04",
  1149 => x"b6b40881",
  1150 => x"e02e0981",
  1151 => x"06893881",
  1152 => x"0bb6ac0c",
  1153 => x"a4dc04b6",
  1154 => x"b40852b6",
  1155 => x"ac08802e",
  1156 => x"8838b6b4",
  1157 => x"08818005",
  1158 => x"5271842c",
  1159 => x"728f0653",
  1160 => x"53b6a808",
  1161 => x"802e9938",
  1162 => x"728429b5",
  1163 => x"e8057213",
  1164 => x"81712b70",
  1165 => x"09730806",
  1166 => x"730c5153",
  1167 => x"53a4d204",
  1168 => x"728429b5",
  1169 => x"e8057213",
  1170 => x"83712b72",
  1171 => x"0807720c",
  1172 => x"5353800b",
  1173 => x"b6ac0c80",
  1174 => x"0bb6a80c",
  1175 => x"bce851a2",
  1176 => x"a02db6b4",
  1177 => x"08ff24fe",
  1178 => x"f838800b",
  1179 => x"b6b40c02",
  1180 => x"8c050d04",
  1181 => x"02f8050d",
  1182 => x"b5e8528f",
  1183 => x"51807270",
  1184 => x"8405540c",
  1185 => x"ff115170",
  1186 => x"8025f238",
  1187 => x"0288050d",
  1188 => x"0402f005",
  1189 => x"0d7551a5",
  1190 => x"db2d7082",
  1191 => x"2cfc06b5",
  1192 => x"e8117210",
  1193 => x"9e067108",
  1194 => x"70722a70",
  1195 => x"83068274",
  1196 => x"2b700974",
  1197 => x"06760c54",
  1198 => x"51565753",
  1199 => x"5153a5d5",
  1200 => x"2d71b6b4",
  1201 => x"0c029005",
  1202 => x"0d047198",
  1203 => x"0c04ffb0",
  1204 => x"08b6b40c",
  1205 => x"04810bff",
  1206 => x"b00c0480",
  1207 => x"0bffb00c",
  1208 => x"0402fc05",
  1209 => x"0d810bb6",
  1210 => x"b00c8151",
  1211 => x"84e52d02",
  1212 => x"84050d04",
  1213 => x"02fc050d",
  1214 => x"800bb6b0",
  1215 => x"0c805184",
  1216 => x"e52d0284",
  1217 => x"050d0402",
  1218 => x"ec050d76",
  1219 => x"54805287",
  1220 => x"0b881580",
  1221 => x"f52d5653",
  1222 => x"74722483",
  1223 => x"38a05372",
  1224 => x"5182ee2d",
  1225 => x"81128b15",
  1226 => x"80f52d54",
  1227 => x"52727225",
  1228 => x"de380294",
  1229 => x"050d0402",
  1230 => x"f0050dbd",
  1231 => x"a0085481",
  1232 => x"f72d800b",
  1233 => x"bda40c73",
  1234 => x"08802e81",
  1235 => x"8038820b",
  1236 => x"b6c80cbd",
  1237 => x"a4088f06",
  1238 => x"b6c40c73",
  1239 => x"08527183",
  1240 => x"2e963871",
  1241 => x"83268938",
  1242 => x"71812eaf",
  1243 => x"38a7b804",
  1244 => x"71852e9f",
  1245 => x"38a7b804",
  1246 => x"881480f5",
  1247 => x"2d841508",
  1248 => x"b3985354",
  1249 => x"5285f12d",
  1250 => x"71842913",
  1251 => x"70085252",
  1252 => x"a7bc0473",
  1253 => x"51a6872d",
  1254 => x"a7b804bd",
  1255 => x"94088815",
  1256 => x"082c7081",
  1257 => x"06515271",
  1258 => x"802e8738",
  1259 => x"b39c51a7",
  1260 => x"b504b3a0",
  1261 => x"5185f12d",
  1262 => x"84140851",
  1263 => x"85f12dbd",
  1264 => x"a4088105",
  1265 => x"bda40c8c",
  1266 => x"1454a6c7",
  1267 => x"04029005",
  1268 => x"0d0471bd",
  1269 => x"a00ca6b7",
  1270 => x"2dbda408",
  1271 => x"ff05bda8",
  1272 => x"0c0471bd",
  1273 => x"ac0c0402",
  1274 => x"e8050dbd",
  1275 => x"a008bdac",
  1276 => x"08575580",
  1277 => x"f851a591",
  1278 => x"2db6b408",
  1279 => x"812a7081",
  1280 => x"06515271",
  1281 => x"9b388751",
  1282 => x"a5912db6",
  1283 => x"b408812a",
  1284 => x"70810651",
  1285 => x"5271802e",
  1286 => x"b138a8a0",
  1287 => x"04a3da2d",
  1288 => x"8751a591",
  1289 => x"2db6b408",
  1290 => x"f438a8b0",
  1291 => x"04a3da2d",
  1292 => x"80f851a5",
  1293 => x"912db6b4",
  1294 => x"08f338b6",
  1295 => x"b0088132",
  1296 => x"70b6b00c",
  1297 => x"70525284",
  1298 => x"e52d800b",
  1299 => x"bd980c80",
  1300 => x"0bbd9c0c",
  1301 => x"b6b00882",
  1302 => x"dd3880da",
  1303 => x"51a5912d",
  1304 => x"b6b40880",
  1305 => x"2e8a38bd",
  1306 => x"98088180",
  1307 => x"07bd980c",
  1308 => x"80d951a5",
  1309 => x"912db6b4",
  1310 => x"08802e8a",
  1311 => x"38bd9808",
  1312 => x"80c007bd",
  1313 => x"980c8194",
  1314 => x"51a5912d",
  1315 => x"b6b40880",
  1316 => x"2e8938bd",
  1317 => x"98089007",
  1318 => x"bd980c81",
  1319 => x"9151a591",
  1320 => x"2db6b408",
  1321 => x"802e8938",
  1322 => x"bd9808a0",
  1323 => x"07bd980c",
  1324 => x"81f551a5",
  1325 => x"912db6b4",
  1326 => x"08802e89",
  1327 => x"38bd9808",
  1328 => x"8107bd98",
  1329 => x"0c81f251",
  1330 => x"a5912db6",
  1331 => x"b408802e",
  1332 => x"8938bd98",
  1333 => x"088207bd",
  1334 => x"980c81eb",
  1335 => x"51a5912d",
  1336 => x"b6b40880",
  1337 => x"2e8938bd",
  1338 => x"98088407",
  1339 => x"bd980c81",
  1340 => x"f451a591",
  1341 => x"2db6b408",
  1342 => x"802e8938",
  1343 => x"bd980888",
  1344 => x"07bd980c",
  1345 => x"80d851a5",
  1346 => x"912db6b4",
  1347 => x"08802e8a",
  1348 => x"38bd9c08",
  1349 => x"818007bd",
  1350 => x"9c0c9251",
  1351 => x"a5912db6",
  1352 => x"b408802e",
  1353 => x"8a38bd9c",
  1354 => x"0880c007",
  1355 => x"bd9c0c94",
  1356 => x"51a5912d",
  1357 => x"b6b40880",
  1358 => x"2e8938bd",
  1359 => x"9c089007",
  1360 => x"bd9c0c91",
  1361 => x"51a5912d",
  1362 => x"b6b40880",
  1363 => x"2e8938bd",
  1364 => x"9c08a007",
  1365 => x"bd9c0c9d",
  1366 => x"51a5912d",
  1367 => x"b6b40880",
  1368 => x"2e8938bd",
  1369 => x"9c088107",
  1370 => x"bd9c0c9b",
  1371 => x"51a5912d",
  1372 => x"b6b40880",
  1373 => x"2e8938bd",
  1374 => x"9c088207",
  1375 => x"bd9c0c9c",
  1376 => x"51a5912d",
  1377 => x"b6b40880",
  1378 => x"2e8938bd",
  1379 => x"9c088407",
  1380 => x"bd9c0ca3",
  1381 => x"51a5912d",
  1382 => x"b6b40880",
  1383 => x"2e8938bd",
  1384 => x"9c088807",
  1385 => x"bd9c0c81",
  1386 => x"fd51a591",
  1387 => x"2d81fa51",
  1388 => x"a5912db0",
  1389 => x"9b0481f5",
  1390 => x"51a5912d",
  1391 => x"b6b40881",
  1392 => x"2a708106",
  1393 => x"51527180",
  1394 => x"2eaf38bd",
  1395 => x"a8085271",
  1396 => x"802e8938",
  1397 => x"ff12bda8",
  1398 => x"0cabf904",
  1399 => x"bda40810",
  1400 => x"bda40805",
  1401 => x"70842916",
  1402 => x"51528812",
  1403 => x"08802e89",
  1404 => x"38ff5188",
  1405 => x"12085271",
  1406 => x"2d81f251",
  1407 => x"a5912db6",
  1408 => x"b408812a",
  1409 => x"70810651",
  1410 => x"5271802e",
  1411 => x"b138bda4",
  1412 => x"08ff11bd",
  1413 => x"a8085653",
  1414 => x"53737225",
  1415 => x"89388114",
  1416 => x"bda80cac",
  1417 => x"be047210",
  1418 => x"13708429",
  1419 => x"16515288",
  1420 => x"1208802e",
  1421 => x"8938fe51",
  1422 => x"88120852",
  1423 => x"712d81fd",
  1424 => x"51a5912d",
  1425 => x"b6b40881",
  1426 => x"2a708106",
  1427 => x"51527180",
  1428 => x"2e863880",
  1429 => x"0bbda80c",
  1430 => x"81fa51a5",
  1431 => x"912db6b4",
  1432 => x"08812a70",
  1433 => x"81065152",
  1434 => x"71802e89",
  1435 => x"38bda408",
  1436 => x"ff05bda8",
  1437 => x"0cbda808",
  1438 => x"70535473",
  1439 => x"802e8a38",
  1440 => x"8c15ff15",
  1441 => x"5555acfb",
  1442 => x"04820bb6",
  1443 => x"c80c718f",
  1444 => x"06b6c40c",
  1445 => x"81eb51a5",
  1446 => x"912db6b4",
  1447 => x"08812a70",
  1448 => x"81065152",
  1449 => x"71802ead",
  1450 => x"38740885",
  1451 => x"2e098106",
  1452 => x"a4388815",
  1453 => x"80f52dff",
  1454 => x"05527188",
  1455 => x"1681b72d",
  1456 => x"71982b52",
  1457 => x"71802588",
  1458 => x"38800b88",
  1459 => x"1681b72d",
  1460 => x"7451a687",
  1461 => x"2d81f451",
  1462 => x"a5912db6",
  1463 => x"b408812a",
  1464 => x"70810651",
  1465 => x"5271802e",
  1466 => x"b3387408",
  1467 => x"852e0981",
  1468 => x"06aa3888",
  1469 => x"1580f52d",
  1470 => x"81055271",
  1471 => x"881681b7",
  1472 => x"2d7181ff",
  1473 => x"068b1680",
  1474 => x"f52d5452",
  1475 => x"72722787",
  1476 => x"38728816",
  1477 => x"81b72d74",
  1478 => x"51a6872d",
  1479 => x"80da51a5",
  1480 => x"912db6b4",
  1481 => x"08812a70",
  1482 => x"81065152",
  1483 => x"71802e81",
  1484 => x"a638bda0",
  1485 => x"08bda808",
  1486 => x"55537380",
  1487 => x"2e8a388c",
  1488 => x"13ff1555",
  1489 => x"53aeba04",
  1490 => x"72085271",
  1491 => x"822ea638",
  1492 => x"71822689",
  1493 => x"3871812e",
  1494 => x"a938afd7",
  1495 => x"0471832e",
  1496 => x"b1387184",
  1497 => x"2e098106",
  1498 => x"80ed3888",
  1499 => x"130851a7",
  1500 => x"d22dafd7",
  1501 => x"04bda808",
  1502 => x"51881308",
  1503 => x"52712daf",
  1504 => x"d704810b",
  1505 => x"8814082b",
  1506 => x"bd940832",
  1507 => x"bd940caf",
  1508 => x"ad048813",
  1509 => x"80f52d81",
  1510 => x"058b1480",
  1511 => x"f52d5354",
  1512 => x"71742483",
  1513 => x"38805473",
  1514 => x"881481b7",
  1515 => x"2da6b72d",
  1516 => x"afd70475",
  1517 => x"08802ea2",
  1518 => x"38750851",
  1519 => x"a5912db6",
  1520 => x"b4088106",
  1521 => x"5271802e",
  1522 => x"8b38bda8",
  1523 => x"08518416",
  1524 => x"0852712d",
  1525 => x"88165675",
  1526 => x"da388054",
  1527 => x"800bb6c8",
  1528 => x"0c738f06",
  1529 => x"b6c40ca0",
  1530 => x"5273bda8",
  1531 => x"082e0981",
  1532 => x"069838bd",
  1533 => x"a408ff05",
  1534 => x"74327009",
  1535 => x"81057072",
  1536 => x"079f2a91",
  1537 => x"71315151",
  1538 => x"53537151",
  1539 => x"82ee2d81",
  1540 => x"14548e74",
  1541 => x"25c638b6",
  1542 => x"b0085271",
  1543 => x"b6b40c02",
  1544 => x"98050d04",
  1545 => x"00ffffff",
  1546 => x"ff00ffff",
  1547 => x"ffff00ff",
  1548 => x"ffffff00",
  1549 => x"52657365",
  1550 => x"74000000",
  1551 => x"53617665",
  1552 => x"20736574",
  1553 => x"74696e67",
  1554 => x"73000000",
  1555 => x"5363616e",
  1556 => x"6c696e65",
  1557 => x"73000000",
  1558 => x"4c6f6164",
  1559 => x"20524f4d",
  1560 => x"20100000",
  1561 => x"45786974",
  1562 => x"00000000",
  1563 => x"50432045",
  1564 => x"6e67696e",
  1565 => x"65206d6f",
  1566 => x"64650000",
  1567 => x"54757262",
  1568 => x"6f677261",
  1569 => x"66782031",
  1570 => x"36206d6f",
  1571 => x"64650000",
  1572 => x"56474120",
  1573 => x"2d203331",
  1574 => x"4b487a2c",
  1575 => x"20363048",
  1576 => x"7a000000",
  1577 => x"5456202d",
  1578 => x"20343830",
  1579 => x"692c2036",
  1580 => x"30487a00",
  1581 => x"4261636b",
  1582 => x"00000000",
  1583 => x"46504741",
  1584 => x"50434520",
  1585 => x"43464700",
  1586 => x"496e6974",
  1587 => x"69616c69",
  1588 => x"7a696e67",
  1589 => x"20534420",
  1590 => x"63617264",
  1591 => x"0a000000",
  1592 => x"424f4f54",
  1593 => x"20202020",
  1594 => x"50434500",
  1595 => x"43617264",
  1596 => x"20696e69",
  1597 => x"74206661",
  1598 => x"696c6564",
  1599 => x"0a000000",
  1600 => x"4d425220",
  1601 => x"6661696c",
  1602 => x"0a000000",
  1603 => x"46415431",
  1604 => x"36202020",
  1605 => x"00000000",
  1606 => x"46415433",
  1607 => x"32202020",
  1608 => x"00000000",
  1609 => x"4e6f2070",
  1610 => x"61727469",
  1611 => x"74696f6e",
  1612 => x"20736967",
  1613 => x"0a000000",
  1614 => x"42616420",
  1615 => x"70617274",
  1616 => x"0a000000",
  1617 => x"53444843",
  1618 => x"20657272",
  1619 => x"6f72210a",
  1620 => x"00000000",
  1621 => x"53442069",
  1622 => x"6e69742e",
  1623 => x"2e2e0a00",
  1624 => x"53442063",
  1625 => x"61726420",
  1626 => x"72657365",
  1627 => x"74206661",
  1628 => x"696c6564",
  1629 => x"210a0000",
  1630 => x"57726974",
  1631 => x"65206661",
  1632 => x"696c6564",
  1633 => x"0a000000",
  1634 => x"52656164",
  1635 => x"20666169",
  1636 => x"6c65640a",
  1637 => x"00000000",
  1638 => x"16200000",
  1639 => x"14200000",
  1640 => x"15200000",
  1641 => x"00000002",
  1642 => x"00000002",
  1643 => x"00001834",
  1644 => x"000004b0",
  1645 => x"00000002",
  1646 => x"0000183c",
  1647 => x"00000377",
  1648 => x"00000003",
  1649 => x"00001a10",
  1650 => x"00000002",
  1651 => x"00000001",
  1652 => x"0000184c",
  1653 => x"00000001",
  1654 => x"00000003",
  1655 => x"00001a08",
  1656 => x"00000002",
  1657 => x"00000002",
  1658 => x"00001858",
  1659 => x"00000631",
  1660 => x"00000002",
  1661 => x"00001864",
  1662 => x"000012f4",
  1663 => x"00000000",
  1664 => x"00000000",
  1665 => x"00000000",
  1666 => x"0000186c",
  1667 => x"0000187c",
  1668 => x"00001890",
  1669 => x"000018a4",
  1670 => x"0000004d",
  1671 => x"00000605",
  1672 => x"0000002c",
  1673 => x"0000061b",
  1674 => x"00000000",
  1675 => x"00000000",
  1676 => x"00000002",
  1677 => x"00001b64",
  1678 => x"000004c5",
  1679 => x"00000002",
  1680 => x"00001b74",
  1681 => x"000004c5",
  1682 => x"00000002",
  1683 => x"00001b84",
  1684 => x"000004c5",
  1685 => x"00000002",
  1686 => x"00001b94",
  1687 => x"000004c5",
  1688 => x"00000002",
  1689 => x"00001ba4",
  1690 => x"000004c5",
  1691 => x"00000002",
  1692 => x"00001bb4",
  1693 => x"000004c5",
  1694 => x"00000002",
  1695 => x"00001bc4",
  1696 => x"000004c5",
  1697 => x"00000002",
  1698 => x"00001bd4",
  1699 => x"000004c5",
  1700 => x"00000002",
  1701 => x"00001be4",
  1702 => x"000004c5",
  1703 => x"00000002",
  1704 => x"00001bf4",
  1705 => x"000004c5",
  1706 => x"00000002",
  1707 => x"00001c04",
  1708 => x"000004c5",
  1709 => x"00000002",
  1710 => x"00001c14",
  1711 => x"000004c5",
  1712 => x"00000002",
  1713 => x"00001c24",
  1714 => x"000004c5",
  1715 => x"00000004",
  1716 => x"000018b4",
  1717 => x"000019a8",
  1718 => x"00000000",
  1719 => x"00000000",
  1720 => x"00000599",
  1721 => x"00000000",
  1722 => x"00000000",
  1723 => x"00000000",
  1724 => x"00000000",
  1725 => x"00000000",
  1726 => x"00000000",
  1727 => x"00000000",
  1728 => x"00000000",
  1729 => x"00000000",
  1730 => x"00000000",
  1731 => x"00000000",
  1732 => x"00000000",
  1733 => x"00000000",
  1734 => x"00000000",
  1735 => x"00000000",
  1736 => x"00000000",
  1737 => x"00000000",
  1738 => x"00000000",
  1739 => x"00000000",
  1740 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

