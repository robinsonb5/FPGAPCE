-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb5",
     9 => x"d8080b0b",
    10 => x"0bb5dc08",
    11 => x"0b0b0bb5",
    12 => x"e0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b5e00c0b",
    16 => x"0b0bb5dc",
    17 => x"0c0b0b0b",
    18 => x"b5d80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bafcc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b5d870bc",
    57 => x"d4278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8ce20402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b5e80c9f",
    65 => x"0bb5ec0c",
    66 => x"a0717081",
    67 => x"055334b5",
    68 => x"ec08ff05",
    69 => x"b5ec0cb5",
    70 => x"ec088025",
    71 => x"eb38b5e8",
    72 => x"08ff05b5",
    73 => x"e80cb5e8",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb5e8",
    94 => x"08258f38",
    95 => x"82b22db5",
    96 => x"e808ff05",
    97 => x"b5e80c82",
    98 => x"f404b5e8",
    99 => x"08b5ec08",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b5e808",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b5",
   108 => x"ec088105",
   109 => x"b5ec0cb5",
   110 => x"ec08519f",
   111 => x"7125e238",
   112 => x"800bb5ec",
   113 => x"0cb5e808",
   114 => x"8105b5e8",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b5ec0881",
   120 => x"05b5ec0c",
   121 => x"b5ec08a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b5ec0cb5",
   125 => x"e8088105",
   126 => x"b5e80c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb5",
   155 => x"f00cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb5f0",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b5f00884",
   167 => x"07b5f00c",
   168 => x"5573842b",
   169 => x"87e87125",
   170 => x"83713170",
   171 => x"0b0b0bb2",
   172 => x"e00c8171",
   173 => x"2bf6880c",
   174 => x"fea413ff",
   175 => x"122c7888",
   176 => x"29ff9405",
   177 => x"70812cb5",
   178 => x"f0085258",
   179 => x"52555152",
   180 => x"5476802e",
   181 => x"85387081",
   182 => x"075170f6",
   183 => x"940c7109",
   184 => x"8105f680",
   185 => x"0c720981",
   186 => x"05f6840c",
   187 => x"0294050d",
   188 => x"0402f405",
   189 => x"0d745372",
   190 => x"70810554",
   191 => x"80f52d52",
   192 => x"71802e89",
   193 => x"38715182",
   194 => x"ee2d85f7",
   195 => x"04028c05",
   196 => x"0d0402f4",
   197 => x"050d7470",
   198 => x"8206bcbc",
   199 => x"0cb2fc71",
   200 => x"81065454",
   201 => x"51718814",
   202 => x"81b72d70",
   203 => x"822a7081",
   204 => x"06515170",
   205 => x"941481b7",
   206 => x"2d70b5d8",
   207 => x"0c028c05",
   208 => x"0d0402f4",
   209 => x"050db0e4",
   210 => x"52b5f851",
   211 => x"96852db5",
   212 => x"d808802e",
   213 => x"9538b7dc",
   214 => x"52b5f851",
   215 => x"98bb2db7",
   216 => x"dc0870fe",
   217 => x"c00c5186",
   218 => x"922d028c",
   219 => x"050d0402",
   220 => x"f8050dbc",
   221 => x"bc088206",
   222 => x"b3840b80",
   223 => x"f52d5252",
   224 => x"70802e85",
   225 => x"38718107",
   226 => x"52b39c0b",
   227 => x"80f52d51",
   228 => x"70802e85",
   229 => x"38718407",
   230 => x"5271b684",
   231 => x"080752b6",
   232 => x"8808802e",
   233 => x"85387190",
   234 => x"075271b5",
   235 => x"d80c0288",
   236 => x"050d0402",
   237 => x"f0050d86",
   238 => x"ef2db5d8",
   239 => x"08b0e453",
   240 => x"b5f85253",
   241 => x"96852db5",
   242 => x"d808802e",
   243 => x"a33872b7",
   244 => x"dc0cb7e0",
   245 => x"5480fd53",
   246 => x"80747084",
   247 => x"05560cff",
   248 => x"13537280",
   249 => x"25f238b7",
   250 => x"dc52b5f8",
   251 => x"5198e12d",
   252 => x"0290050d",
   253 => x"0402d805",
   254 => x"0d810bfe",
   255 => x"c40c840b",
   256 => x"fec40c7b",
   257 => x"52b5f851",
   258 => x"96852db5",
   259 => x"d80853b5",
   260 => x"d808802e",
   261 => x"81c638b5",
   262 => x"fc085680",
   263 => x"0bff1758",
   264 => x"5976792e",
   265 => x"8b388119",
   266 => x"77812a58",
   267 => x"5976f738",
   268 => x"f719769f",
   269 => x"ff065459",
   270 => x"72802e8b",
   271 => x"38fc8016",
   272 => x"b5f85256",
   273 => x"988e2d75",
   274 => x"b080802e",
   275 => x"09810689",
   276 => x"38880bb6",
   277 => x"840c88e6",
   278 => x"04800bb6",
   279 => x"840c8153",
   280 => x"80762580",
   281 => x"fd387852",
   282 => x"76518480",
   283 => x"2db7dc52",
   284 => x"b5f85198",
   285 => x"bb2db5d8",
   286 => x"08b7dc5b",
   287 => x"538058b5",
   288 => x"d808b038",
   289 => x"89c60479",
   290 => x"7084055b",
   291 => x"087083fe",
   292 => x"80067188",
   293 => x"2b83fe80",
   294 => x"0671882a",
   295 => x"0772882a",
   296 => x"83fe8006",
   297 => x"73982a07",
   298 => x"fec80cfe",
   299 => x"c80c5684",
   300 => x"19595375",
   301 => x"53848076",
   302 => x"25843884",
   303 => x"80537278",
   304 => x"24c53889",
   305 => x"cc04b0f0",
   306 => x"5189df04",
   307 => x"b5f85198",
   308 => x"8e2dfc80",
   309 => x"16811858",
   310 => x"5688de04",
   311 => x"b1805185",
   312 => x"f12d72b5",
   313 => x"d80c02a8",
   314 => x"050d0402",
   315 => x"fc050da5",
   316 => x"cf2dfec4",
   317 => x"5181710c",
   318 => x"82710c02",
   319 => x"84050d04",
   320 => x"02f4050d",
   321 => x"74101570",
   322 => x"8429b3d8",
   323 => x"05700855",
   324 => x"51527280",
   325 => x"2e9b3872",
   326 => x"80f52d52",
   327 => x"71802e91",
   328 => x"38b18851",
   329 => x"85f12d72",
   330 => x"5185f12d",
   331 => x"725187f5",
   332 => x"2db2e451",
   333 => x"a7ad2da5",
   334 => x"cf2d8051",
   335 => x"84e52d02",
   336 => x"8c050d04",
   337 => x"02e8050d",
   338 => x"80705656",
   339 => x"75b58808",
   340 => x"25af38bb",
   341 => x"e808762e",
   342 => x"a8387451",
   343 => x"95b02db5",
   344 => x"d8080981",
   345 => x"0570b5d8",
   346 => x"08079f2a",
   347 => x"77058117",
   348 => x"57575275",
   349 => x"b5880825",
   350 => x"8838bbe8",
   351 => x"087526da",
   352 => x"38805674",
   353 => x"bbe80827",
   354 => x"80d03874",
   355 => x"5195b02d",
   356 => x"75842b52",
   357 => x"b5d80880",
   358 => x"2eae38b6",
   359 => x"8c128117",
   360 => x"b5d80856",
   361 => x"57528a53",
   362 => x"73708105",
   363 => x"5580f52d",
   364 => x"72708105",
   365 => x"5481b72d",
   366 => x"ff135372",
   367 => x"8025e938",
   368 => x"807281b7",
   369 => x"2d8bd104",
   370 => x"b5d808b6",
   371 => x"8c1381b7",
   372 => x"2d811555",
   373 => x"8b7625ff",
   374 => x"aa380298",
   375 => x"050d0402",
   376 => x"fc050d72",
   377 => x"5170fd2e",
   378 => x"ad3870fd",
   379 => x"248a3870",
   380 => x"fc2e80c4",
   381 => x"388cc004",
   382 => x"70fe2eb1",
   383 => x"3870ff2e",
   384 => x"098106bc",
   385 => x"38b58808",
   386 => x"5170802e",
   387 => x"b338ff11",
   388 => x"b5880c8c",
   389 => x"c004b588",
   390 => x"08f00570",
   391 => x"b5880c51",
   392 => x"7080259c",
   393 => x"38800bb5",
   394 => x"880c8cc0",
   395 => x"04b58808",
   396 => x"8105b588",
   397 => x"0c8cc004",
   398 => x"b5880890",
   399 => x"05b5880c",
   400 => x"8ac42da6",
   401 => x"922d0284",
   402 => x"050d0402",
   403 => x"fc050d80",
   404 => x"0bb5880c",
   405 => x"8ac42db3",
   406 => x"d451a7ad",
   407 => x"2d028405",
   408 => x"0d0402f4",
   409 => x"050d800b",
   410 => x"b6840c81",
   411 => x"0bb6880c",
   412 => x"90518692",
   413 => x"2d810bfe",
   414 => x"c40c900b",
   415 => x"fec00c84",
   416 => x"0bfec40c",
   417 => x"830bfecc",
   418 => x"0ca39d2d",
   419 => x"a5b02da3",
   420 => x"822da382",
   421 => x"2d81f72d",
   422 => x"815184e5",
   423 => x"2da3822d",
   424 => x"a3822d81",
   425 => x"5184e52d",
   426 => x"b1945185",
   427 => x"f12d8452",
   428 => x"9d942d8f",
   429 => x"9e2db5d8",
   430 => x"08802e86",
   431 => x"38fe528d",
   432 => x"ca04ff12",
   433 => x"52718024",
   434 => x"e7387180",
   435 => x"2e818138",
   436 => x"86c22db1",
   437 => x"ac5187f5",
   438 => x"2db5d808",
   439 => x"802e8f38",
   440 => x"b2e451a7",
   441 => x"ad2d8051",
   442 => x"84e52d8d",
   443 => x"f804b5d8",
   444 => x"08518ccb",
   445 => x"2da5bc2d",
   446 => x"a3b52da7",
   447 => x"bd2db5d8",
   448 => x"08bcc008",
   449 => x"882bbcc4",
   450 => x"0807fed8",
   451 => x"0c5386ef",
   452 => x"2db5d808",
   453 => x"b5f4082e",
   454 => x"a238b5d8",
   455 => x"08b5f40c",
   456 => x"b5d808fe",
   457 => x"c00c8452",
   458 => x"725184e5",
   459 => x"2da3822d",
   460 => x"a3822dff",
   461 => x"12527180",
   462 => x"25ee3872",
   463 => x"802e8938",
   464 => x"8a0bfec4",
   465 => x"0c8df804",
   466 => x"820bfec4",
   467 => x"0c8df804",
   468 => x"b1b85185",
   469 => x"f12d800b",
   470 => x"b5d80c02",
   471 => x"8c050d04",
   472 => x"02e8050d",
   473 => x"77797b58",
   474 => x"55558053",
   475 => x"727625a3",
   476 => x"38747081",
   477 => x"055680f5",
   478 => x"2d747081",
   479 => x"055680f5",
   480 => x"2d525271",
   481 => x"712e8638",
   482 => x"81518f95",
   483 => x"04811353",
   484 => x"8eec0480",
   485 => x"5170b5d8",
   486 => x"0c029805",
   487 => x"0d0402d8",
   488 => x"050d800b",
   489 => x"bbe40cb7",
   490 => x"dc528051",
   491 => x"9ffc2db5",
   492 => x"d80854b5",
   493 => x"d8088c38",
   494 => x"b1cc5185",
   495 => x"f12d7355",
   496 => x"94b90480",
   497 => x"56810bbc",
   498 => x"880c8853",
   499 => x"b1d852b8",
   500 => x"92518ee0",
   501 => x"2db5d808",
   502 => x"762e0981",
   503 => x"068738b5",
   504 => x"d808bc88",
   505 => x"0c8853b1",
   506 => x"e452b8ae",
   507 => x"518ee02d",
   508 => x"b5d80887",
   509 => x"38b5d808",
   510 => x"bc880cbc",
   511 => x"8808802e",
   512 => x"80f638bb",
   513 => x"a20b80f5",
   514 => x"2dbba30b",
   515 => x"80f52d71",
   516 => x"982b7190",
   517 => x"2b07bba4",
   518 => x"0b80f52d",
   519 => x"70882b72",
   520 => x"07bba50b",
   521 => x"80f52d71",
   522 => x"07bbda0b",
   523 => x"80f52dbb",
   524 => x"db0b80f5",
   525 => x"2d71882b",
   526 => x"07535f54",
   527 => x"525a5657",
   528 => x"557381ab",
   529 => x"aa2e0981",
   530 => x"068d3875",
   531 => x"51a19c2d",
   532 => x"b5d80856",
   533 => x"90e40473",
   534 => x"82d4d52e",
   535 => x"8738b1f0",
   536 => x"5191a504",
   537 => x"b7dc5275",
   538 => x"519ffc2d",
   539 => x"b5d80855",
   540 => x"b5d80880",
   541 => x"2e83c238",
   542 => x"8853b1e4",
   543 => x"52b8ae51",
   544 => x"8ee02db5",
   545 => x"d8088938",
   546 => x"810bbbe4",
   547 => x"0c91ab04",
   548 => x"8853b1d8",
   549 => x"52b89251",
   550 => x"8ee02db5",
   551 => x"d808802e",
   552 => x"8a38b284",
   553 => x"5185f12d",
   554 => x"928504bb",
   555 => x"da0b80f5",
   556 => x"2d547380",
   557 => x"d52e0981",
   558 => x"0680ca38",
   559 => x"bbdb0b80",
   560 => x"f52d5473",
   561 => x"81aa2e09",
   562 => x"8106ba38",
   563 => x"800bb7dc",
   564 => x"0b80f52d",
   565 => x"56547481",
   566 => x"e92e8338",
   567 => x"81547481",
   568 => x"eb2e8c38",
   569 => x"80557375",
   570 => x"2e098106",
   571 => x"82cb38b7",
   572 => x"e70b80f5",
   573 => x"2d55748d",
   574 => x"38b7e80b",
   575 => x"80f52d54",
   576 => x"73822e86",
   577 => x"38805594",
   578 => x"b904b7e9",
   579 => x"0b80f52d",
   580 => x"70bbdc0c",
   581 => x"ff05bbe0",
   582 => x"0cb7ea0b",
   583 => x"80f52db7",
   584 => x"eb0b80f5",
   585 => x"2d587605",
   586 => x"77828029",
   587 => x"0570bbec",
   588 => x"0cb7ec0b",
   589 => x"80f52d70",
   590 => x"bc800cbb",
   591 => x"e4085957",
   592 => x"5876802e",
   593 => x"81a33888",
   594 => x"53b1e452",
   595 => x"b8ae518e",
   596 => x"e02db5d8",
   597 => x"0881e238",
   598 => x"bbdc0870",
   599 => x"842bbbe8",
   600 => x"0c70bbfc",
   601 => x"0cb8810b",
   602 => x"80f52db8",
   603 => x"800b80f5",
   604 => x"2d718280",
   605 => x"2905b882",
   606 => x"0b80f52d",
   607 => x"70848080",
   608 => x"2912b883",
   609 => x"0b80f52d",
   610 => x"7081800a",
   611 => x"291270bc",
   612 => x"840cbc80",
   613 => x"087129bb",
   614 => x"ec080570",
   615 => x"bbf00cb8",
   616 => x"890b80f5",
   617 => x"2db8880b",
   618 => x"80f52d71",
   619 => x"82802905",
   620 => x"b88a0b80",
   621 => x"f52d7084",
   622 => x"80802912",
   623 => x"b88b0b80",
   624 => x"f52d7098",
   625 => x"2b81f00a",
   626 => x"06720570",
   627 => x"bbf40cfe",
   628 => x"117e2977",
   629 => x"05bbf80c",
   630 => x"52595243",
   631 => x"545e5152",
   632 => x"59525d57",
   633 => x"595794b7",
   634 => x"04b7ee0b",
   635 => x"80f52db7",
   636 => x"ed0b80f5",
   637 => x"2d718280",
   638 => x"290570bb",
   639 => x"e80c70a0",
   640 => x"2983ff05",
   641 => x"70892a70",
   642 => x"bbfc0cb7",
   643 => x"f30b80f5",
   644 => x"2db7f20b",
   645 => x"80f52d71",
   646 => x"82802905",
   647 => x"70bc840c",
   648 => x"7b71291e",
   649 => x"70bbf80c",
   650 => x"7dbbf40c",
   651 => x"7305bbf0",
   652 => x"0c555e51",
   653 => x"51555581",
   654 => x"5574b5d8",
   655 => x"0c02a805",
   656 => x"0d0402ec",
   657 => x"050d7670",
   658 => x"872c7180",
   659 => x"ff065556",
   660 => x"54bbe408",
   661 => x"8a387388",
   662 => x"2c7481ff",
   663 => x"065455b7",
   664 => x"dc52bbec",
   665 => x"0815519f",
   666 => x"fc2db5d8",
   667 => x"0854b5d8",
   668 => x"08802eb3",
   669 => x"38bbe408",
   670 => x"802e9838",
   671 => x"728429b7",
   672 => x"dc057008",
   673 => x"5253a19c",
   674 => x"2db5d808",
   675 => x"f00a0653",
   676 => x"95a50472",
   677 => x"10b7dc05",
   678 => x"7080e02d",
   679 => x"5253a1cc",
   680 => x"2db5d808",
   681 => x"53725473",
   682 => x"b5d80c02",
   683 => x"94050d04",
   684 => x"02ec050d",
   685 => x"7670842c",
   686 => x"bbf80805",
   687 => x"718f0652",
   688 => x"55537289",
   689 => x"38b7dc52",
   690 => x"73519ffc",
   691 => x"2d72a029",
   692 => x"b7dc0554",
   693 => x"807480f5",
   694 => x"2d545572",
   695 => x"752e8338",
   696 => x"81557281",
   697 => x"e52e9338",
   698 => x"74802e8e",
   699 => x"388b1480",
   700 => x"f52d9806",
   701 => x"5372802e",
   702 => x"83388054",
   703 => x"73b5d80c",
   704 => x"0294050d",
   705 => x"0402cc05",
   706 => x"0d7e605e",
   707 => x"5a800bbb",
   708 => x"f408bbf8",
   709 => x"08595c56",
   710 => x"8058bbe8",
   711 => x"08782e81",
   712 => x"ae38778f",
   713 => x"06a01757",
   714 => x"54738f38",
   715 => x"b7dc5276",
   716 => x"51811757",
   717 => x"9ffc2db7",
   718 => x"dc568076",
   719 => x"80f52d56",
   720 => x"5474742e",
   721 => x"83388154",
   722 => x"7481e52e",
   723 => x"80f63881",
   724 => x"70750655",
   725 => x"5c73802e",
   726 => x"80ea388b",
   727 => x"1680f52d",
   728 => x"98065978",
   729 => x"80de388b",
   730 => x"537c5275",
   731 => x"518ee02d",
   732 => x"b5d80880",
   733 => x"cf389c16",
   734 => x"0851a19c",
   735 => x"2db5d808",
   736 => x"841b0c9a",
   737 => x"1680e02d",
   738 => x"51a1cc2d",
   739 => x"b5d808b5",
   740 => x"d808881c",
   741 => x"0cb5d808",
   742 => x"5555bbe4",
   743 => x"08802e98",
   744 => x"38941680",
   745 => x"e02d51a1",
   746 => x"cc2db5d8",
   747 => x"08902b83",
   748 => x"fff00a06",
   749 => x"70165154",
   750 => x"73881b0c",
   751 => x"787a0c7b",
   752 => x"54988504",
   753 => x"811858bb",
   754 => x"e8087826",
   755 => x"fed438bb",
   756 => x"e408802e",
   757 => x"ae387a51",
   758 => x"94c22db5",
   759 => x"d808b5d8",
   760 => x"0880ffff",
   761 => x"fff80655",
   762 => x"5b7380ff",
   763 => x"fffff82e",
   764 => x"9238b5d8",
   765 => x"08fe05bb",
   766 => x"dc0829bb",
   767 => x"f0080557",
   768 => x"96980480",
   769 => x"5473b5d8",
   770 => x"0c02b405",
   771 => x"0d0402f4",
   772 => x"050d7470",
   773 => x"08810571",
   774 => x"0c7008bb",
   775 => x"e0080653",
   776 => x"53718e38",
   777 => x"88130851",
   778 => x"94c22db5",
   779 => x"d8088814",
   780 => x"0c810bb5",
   781 => x"d80c028c",
   782 => x"050d0402",
   783 => x"f0050d75",
   784 => x"881108fe",
   785 => x"05bbdc08",
   786 => x"29bbf008",
   787 => x"117208bb",
   788 => x"e0080605",
   789 => x"79555354",
   790 => x"549ffc2d",
   791 => x"0290050d",
   792 => x"0402f005",
   793 => x"0d758811",
   794 => x"08fe05bb",
   795 => x"dc0829bb",
   796 => x"f0081172",
   797 => x"08bbe008",
   798 => x"06057955",
   799 => x"5354549e",
   800 => x"bc2d0290",
   801 => x"050d0402",
   802 => x"f4050dd4",
   803 => x"5281ff72",
   804 => x"0c710853",
   805 => x"81ff720c",
   806 => x"72882b83",
   807 => x"fe800672",
   808 => x"087081ff",
   809 => x"06515253",
   810 => x"81ff720c",
   811 => x"72710788",
   812 => x"2b720870",
   813 => x"81ff0651",
   814 => x"525381ff",
   815 => x"720c7271",
   816 => x"07882b72",
   817 => x"087081ff",
   818 => x"067207b5",
   819 => x"d80c5253",
   820 => x"028c050d",
   821 => x"0402f405",
   822 => x"0d747671",
   823 => x"81ff06d4",
   824 => x"0c5353bc",
   825 => x"8c088538",
   826 => x"71892b52",
   827 => x"71982ad4",
   828 => x"0c71902a",
   829 => x"7081ff06",
   830 => x"d40c5171",
   831 => x"882a7081",
   832 => x"ff06d40c",
   833 => x"517181ff",
   834 => x"06d40c72",
   835 => x"902a7081",
   836 => x"ff06d40c",
   837 => x"51d40870",
   838 => x"81ff0651",
   839 => x"5182b8bf",
   840 => x"527081ff",
   841 => x"2e098106",
   842 => x"943881ff",
   843 => x"0bd40cd4",
   844 => x"087081ff",
   845 => x"06ff1454",
   846 => x"515171e5",
   847 => x"3870b5d8",
   848 => x"0c028c05",
   849 => x"0d0402fc",
   850 => x"050d81c7",
   851 => x"5181ff0b",
   852 => x"d40cff11",
   853 => x"51708025",
   854 => x"f4380284",
   855 => x"050d0402",
   856 => x"f0050d9a",
   857 => x"c62d8fcf",
   858 => x"53805287",
   859 => x"fc80f751",
   860 => x"99d52db5",
   861 => x"d80854b5",
   862 => x"d808812e",
   863 => x"098106a3",
   864 => x"3881ff0b",
   865 => x"d40c820a",
   866 => x"52849c80",
   867 => x"e95199d5",
   868 => x"2db5d808",
   869 => x"8b3881ff",
   870 => x"0bd40c73",
   871 => x"539ba904",
   872 => x"9ac62dff",
   873 => x"135372c1",
   874 => x"3872b5d8",
   875 => x"0c029005",
   876 => x"0d0402f4",
   877 => x"050d81ff",
   878 => x"0bd40c93",
   879 => x"53805287",
   880 => x"fc80c151",
   881 => x"99d52db5",
   882 => x"d8088b38",
   883 => x"81ff0bd4",
   884 => x"0c81539b",
   885 => x"df049ac6",
   886 => x"2dff1353",
   887 => x"72df3872",
   888 => x"b5d80c02",
   889 => x"8c050d04",
   890 => x"02f0050d",
   891 => x"9ac62d83",
   892 => x"aa52849c",
   893 => x"80c85199",
   894 => x"d52db5d8",
   895 => x"08812e09",
   896 => x"81069238",
   897 => x"99872db5",
   898 => x"d80883ff",
   899 => x"ff065372",
   900 => x"83aa2e97",
   901 => x"389bb22d",
   902 => x"9ca60481",
   903 => x"549d8b04",
   904 => x"b2905185",
   905 => x"f12d8054",
   906 => x"9d8b0481",
   907 => x"ff0bd40c",
   908 => x"b1539adf",
   909 => x"2db5d808",
   910 => x"802e80c0",
   911 => x"38805287",
   912 => x"fc80fa51",
   913 => x"99d52db5",
   914 => x"d808b138",
   915 => x"81ff0bd4",
   916 => x"0cd40853",
   917 => x"81ff0bd4",
   918 => x"0c81ff0b",
   919 => x"d40c81ff",
   920 => x"0bd40c81",
   921 => x"ff0bd40c",
   922 => x"72862a70",
   923 => x"8106b5d8",
   924 => x"08565153",
   925 => x"72802e93",
   926 => x"389c9b04",
   927 => x"72822eff",
   928 => x"9f38ff13",
   929 => x"5372ffaa",
   930 => x"38725473",
   931 => x"b5d80c02",
   932 => x"90050d04",
   933 => x"02f0050d",
   934 => x"810bbc8c",
   935 => x"0c8454d0",
   936 => x"08708f2a",
   937 => x"70810651",
   938 => x"515372f3",
   939 => x"3872d00c",
   940 => x"9ac62db2",
   941 => x"a05185f1",
   942 => x"2dd00870",
   943 => x"8f2a7081",
   944 => x"06515153",
   945 => x"72f33881",
   946 => x"0bd00cb1",
   947 => x"53805284",
   948 => x"d480c051",
   949 => x"99d52db5",
   950 => x"d808812e",
   951 => x"a1387282",
   952 => x"2e098106",
   953 => x"8c38b2ac",
   954 => x"5185f12d",
   955 => x"80539eb3",
   956 => x"04ff1353",
   957 => x"72d738ff",
   958 => x"145473ff",
   959 => x"a2389be8",
   960 => x"2db5d808",
   961 => x"bc8c0cb5",
   962 => x"d8088b38",
   963 => x"815287fc",
   964 => x"80d05199",
   965 => x"d52d81ff",
   966 => x"0bd40cd0",
   967 => x"08708f2a",
   968 => x"70810651",
   969 => x"515372f3",
   970 => x"3872d00c",
   971 => x"81ff0bd4",
   972 => x"0c815372",
   973 => x"b5d80c02",
   974 => x"90050d04",
   975 => x"02e8050d",
   976 => x"785681ff",
   977 => x"0bd40cd0",
   978 => x"08708f2a",
   979 => x"70810651",
   980 => x"515372f3",
   981 => x"3882810b",
   982 => x"d00c81ff",
   983 => x"0bd40c77",
   984 => x"5287fc80",
   985 => x"d85199d5",
   986 => x"2db5d808",
   987 => x"802e8c38",
   988 => x"b2c45185",
   989 => x"f12d8153",
   990 => x"9ff30481",
   991 => x"ff0bd40c",
   992 => x"81fe0bd4",
   993 => x"0c80ff55",
   994 => x"75708405",
   995 => x"57087098",
   996 => x"2ad40c70",
   997 => x"902c7081",
   998 => x"ff06d40c",
   999 => x"5470882c",
  1000 => x"7081ff06",
  1001 => x"d40c5470",
  1002 => x"81ff06d4",
  1003 => x"0c54ff15",
  1004 => x"55748025",
  1005 => x"d33881ff",
  1006 => x"0bd40c81",
  1007 => x"ff0bd40c",
  1008 => x"81ff0bd4",
  1009 => x"0c868da0",
  1010 => x"5481ff0b",
  1011 => x"d40cd408",
  1012 => x"81ff0655",
  1013 => x"748738ff",
  1014 => x"145473ed",
  1015 => x"3881ff0b",
  1016 => x"d40cd008",
  1017 => x"708f2a70",
  1018 => x"81065151",
  1019 => x"5372f338",
  1020 => x"72d00c72",
  1021 => x"b5d80c02",
  1022 => x"98050d04",
  1023 => x"02e8050d",
  1024 => x"78558056",
  1025 => x"81ff0bd4",
  1026 => x"0cd00870",
  1027 => x"8f2a7081",
  1028 => x"06515153",
  1029 => x"72f33882",
  1030 => x"810bd00c",
  1031 => x"81ff0bd4",
  1032 => x"0c775287",
  1033 => x"fc80d151",
  1034 => x"99d52d80",
  1035 => x"dbc6df54",
  1036 => x"b5d80880",
  1037 => x"2e8a38b0",
  1038 => x"f05185f1",
  1039 => x"2da19304",
  1040 => x"81ff0bd4",
  1041 => x"0cd40870",
  1042 => x"81ff0651",
  1043 => x"537281fe",
  1044 => x"2e098106",
  1045 => x"9d3880ff",
  1046 => x"5399872d",
  1047 => x"b5d80875",
  1048 => x"70840557",
  1049 => x"0cff1353",
  1050 => x"728025ed",
  1051 => x"388156a0",
  1052 => x"f804ff14",
  1053 => x"5473c938",
  1054 => x"81ff0bd4",
  1055 => x"0c81ff0b",
  1056 => x"d40cd008",
  1057 => x"708f2a70",
  1058 => x"81065151",
  1059 => x"5372f338",
  1060 => x"72d00c75",
  1061 => x"b5d80c02",
  1062 => x"98050d04",
  1063 => x"02f4050d",
  1064 => x"7470882a",
  1065 => x"83fe8006",
  1066 => x"7072982a",
  1067 => x"0772882b",
  1068 => x"87fc8080",
  1069 => x"0673982b",
  1070 => x"81f00a06",
  1071 => x"71730707",
  1072 => x"b5d80c56",
  1073 => x"51535102",
  1074 => x"8c050d04",
  1075 => x"02f8050d",
  1076 => x"028e0580",
  1077 => x"f52d7488",
  1078 => x"2b077083",
  1079 => x"ffff06b5",
  1080 => x"d80c5102",
  1081 => x"88050d04",
  1082 => x"02fc050d",
  1083 => x"72518071",
  1084 => x"0c800b84",
  1085 => x"120c0284",
  1086 => x"050d0402",
  1087 => x"f0050d75",
  1088 => x"70088412",
  1089 => x"08535353",
  1090 => x"ff547171",
  1091 => x"2ea838a5",
  1092 => x"b62d8413",
  1093 => x"08708429",
  1094 => x"14881170",
  1095 => x"087081ff",
  1096 => x"06841808",
  1097 => x"81118706",
  1098 => x"841a0c53",
  1099 => x"51555151",
  1100 => x"51a5b02d",
  1101 => x"715473b5",
  1102 => x"d80c0290",
  1103 => x"050d0402",
  1104 => x"f8050da5",
  1105 => x"b62de008",
  1106 => x"708b2a70",
  1107 => x"81065152",
  1108 => x"5270802e",
  1109 => x"9d38bc90",
  1110 => x"08708429",
  1111 => x"bc980573",
  1112 => x"81ff0671",
  1113 => x"0c5151bc",
  1114 => x"90088111",
  1115 => x"8706bc90",
  1116 => x"0c51800b",
  1117 => x"bcb80ca5",
  1118 => x"a92da5b0",
  1119 => x"2d028805",
  1120 => x"0d0402fc",
  1121 => x"050da5b6",
  1122 => x"2d810bbc",
  1123 => x"b80ca5b0",
  1124 => x"2dbcb808",
  1125 => x"5170fa38",
  1126 => x"0284050d",
  1127 => x"0402fc05",
  1128 => x"0dbc9051",
  1129 => x"a1e82da2",
  1130 => x"bf51a5a5",
  1131 => x"2da4cf2d",
  1132 => x"0284050d",
  1133 => x"0402f405",
  1134 => x"0da4b704",
  1135 => x"b5d80881",
  1136 => x"f02e0981",
  1137 => x"06893881",
  1138 => x"0bb5cc0c",
  1139 => x"a4b704b5",
  1140 => x"d80881e0",
  1141 => x"2e098106",
  1142 => x"8938810b",
  1143 => x"b5d00ca4",
  1144 => x"b704b5d8",
  1145 => x"0852b5d0",
  1146 => x"08802e88",
  1147 => x"38b5d808",
  1148 => x"81800552",
  1149 => x"71842c72",
  1150 => x"8f065353",
  1151 => x"b5cc0880",
  1152 => x"2e993872",
  1153 => x"8429b58c",
  1154 => x"05721381",
  1155 => x"712b7009",
  1156 => x"73080673",
  1157 => x"0c515353",
  1158 => x"a4ad0472",
  1159 => x"8429b58c",
  1160 => x"05721383",
  1161 => x"712b7208",
  1162 => x"07720c53",
  1163 => x"53800bb5",
  1164 => x"d00c800b",
  1165 => x"b5cc0cbc",
  1166 => x"9051a1fb",
  1167 => x"2db5d808",
  1168 => x"ff24fef8",
  1169 => x"38800bb5",
  1170 => x"d80c028c",
  1171 => x"050d0402",
  1172 => x"f8050db5",
  1173 => x"8c528f51",
  1174 => x"80727084",
  1175 => x"05540cff",
  1176 => x"11517080",
  1177 => x"25f23802",
  1178 => x"88050d04",
  1179 => x"02f0050d",
  1180 => x"7551a5b6",
  1181 => x"2d70822c",
  1182 => x"fc06b58c",
  1183 => x"1172109e",
  1184 => x"06710870",
  1185 => x"722a7083",
  1186 => x"0682742b",
  1187 => x"70097406",
  1188 => x"760c5451",
  1189 => x"56575351",
  1190 => x"53a5b02d",
  1191 => x"71b5d80c",
  1192 => x"0290050d",
  1193 => x"0471980c",
  1194 => x"04ffb008",
  1195 => x"b5d80c04",
  1196 => x"810bffb0",
  1197 => x"0c04800b",
  1198 => x"ffb00c04",
  1199 => x"02fc050d",
  1200 => x"810bb5d4",
  1201 => x"0c815184",
  1202 => x"e52d0284",
  1203 => x"050d0402",
  1204 => x"fc050d80",
  1205 => x"0bb5d40c",
  1206 => x"805184e5",
  1207 => x"2d028405",
  1208 => x"0d0402ec",
  1209 => x"050d7654",
  1210 => x"8052870b",
  1211 => x"881580f5",
  1212 => x"2d565374",
  1213 => x"72248338",
  1214 => x"a0537251",
  1215 => x"82ee2d81",
  1216 => x"128b1580",
  1217 => x"f52d5452",
  1218 => x"727225de",
  1219 => x"38029405",
  1220 => x"0d0402f0",
  1221 => x"050dbcc8",
  1222 => x"085481f7",
  1223 => x"2d800bbc",
  1224 => x"cc0c7308",
  1225 => x"802e8180",
  1226 => x"38820bb5",
  1227 => x"ec0cbccc",
  1228 => x"088f06b5",
  1229 => x"e80c7308",
  1230 => x"5271832e",
  1231 => x"96387183",
  1232 => x"26893871",
  1233 => x"812eaf38",
  1234 => x"a7930471",
  1235 => x"852e9f38",
  1236 => x"a7930488",
  1237 => x"1480f52d",
  1238 => x"841508b2",
  1239 => x"d4535452",
  1240 => x"85f12d71",
  1241 => x"84291370",
  1242 => x"085252a7",
  1243 => x"97047351",
  1244 => x"a5e22da7",
  1245 => x"9304bcbc",
  1246 => x"08881508",
  1247 => x"2c708106",
  1248 => x"51527180",
  1249 => x"2e8738b2",
  1250 => x"d851a790",
  1251 => x"04b2dc51",
  1252 => x"85f12d84",
  1253 => x"14085185",
  1254 => x"f12dbccc",
  1255 => x"088105bc",
  1256 => x"cc0c8c14",
  1257 => x"54a6a204",
  1258 => x"0290050d",
  1259 => x"0471bcc8",
  1260 => x"0ca6922d",
  1261 => x"bccc08ff",
  1262 => x"05bcd00c",
  1263 => x"0402ec05",
  1264 => x"0dbcc808",
  1265 => x"5580f851",
  1266 => x"a4ec2db5",
  1267 => x"d808812a",
  1268 => x"70810651",
  1269 => x"52719b38",
  1270 => x"8751a4ec",
  1271 => x"2db5d808",
  1272 => x"812a7081",
  1273 => x"06515271",
  1274 => x"802eb138",
  1275 => x"a7f204a3",
  1276 => x"b52d8751",
  1277 => x"a4ec2db5",
  1278 => x"d808f438",
  1279 => x"a88204a3",
  1280 => x"b52d80f8",
  1281 => x"51a4ec2d",
  1282 => x"b5d808f3",
  1283 => x"38b5d408",
  1284 => x"813270b5",
  1285 => x"d40c7052",
  1286 => x"5284e52d",
  1287 => x"800bbcc0",
  1288 => x"0c800bbc",
  1289 => x"c40cb5d4",
  1290 => x"0882dd38",
  1291 => x"80da51a4",
  1292 => x"ec2db5d8",
  1293 => x"08802e8a",
  1294 => x"38bcc008",
  1295 => x"818007bc",
  1296 => x"c00c80d9",
  1297 => x"51a4ec2d",
  1298 => x"b5d80880",
  1299 => x"2e8a38bc",
  1300 => x"c00880c0",
  1301 => x"07bcc00c",
  1302 => x"819451a4",
  1303 => x"ec2db5d8",
  1304 => x"08802e89",
  1305 => x"38bcc008",
  1306 => x"9007bcc0",
  1307 => x"0c819151",
  1308 => x"a4ec2db5",
  1309 => x"d808802e",
  1310 => x"8938bcc0",
  1311 => x"08a007bc",
  1312 => x"c00c81f5",
  1313 => x"51a4ec2d",
  1314 => x"b5d80880",
  1315 => x"2e8938bc",
  1316 => x"c0088107",
  1317 => x"bcc00c81",
  1318 => x"f251a4ec",
  1319 => x"2db5d808",
  1320 => x"802e8938",
  1321 => x"bcc00882",
  1322 => x"07bcc00c",
  1323 => x"81eb51a4",
  1324 => x"ec2db5d8",
  1325 => x"08802e89",
  1326 => x"38bcc008",
  1327 => x"8407bcc0",
  1328 => x"0c81f451",
  1329 => x"a4ec2db5",
  1330 => x"d808802e",
  1331 => x"8938bcc0",
  1332 => x"088807bc",
  1333 => x"c00c80d8",
  1334 => x"51a4ec2d",
  1335 => x"b5d80880",
  1336 => x"2e8a38bc",
  1337 => x"c4088180",
  1338 => x"07bcc40c",
  1339 => x"9251a4ec",
  1340 => x"2db5d808",
  1341 => x"802e8a38",
  1342 => x"bcc40880",
  1343 => x"c007bcc4",
  1344 => x"0c9451a4",
  1345 => x"ec2db5d8",
  1346 => x"08802e89",
  1347 => x"38bcc408",
  1348 => x"9007bcc4",
  1349 => x"0c9151a4",
  1350 => x"ec2db5d8",
  1351 => x"08802e89",
  1352 => x"38bcc408",
  1353 => x"a007bcc4",
  1354 => x"0c9d51a4",
  1355 => x"ec2db5d8",
  1356 => x"08802e89",
  1357 => x"38bcc408",
  1358 => x"8107bcc4",
  1359 => x"0c9b51a4",
  1360 => x"ec2db5d8",
  1361 => x"08802e89",
  1362 => x"38bcc408",
  1363 => x"8207bcc4",
  1364 => x"0c9c51a4",
  1365 => x"ec2db5d8",
  1366 => x"08802e89",
  1367 => x"38bcc408",
  1368 => x"8407bcc4",
  1369 => x"0ca351a4",
  1370 => x"ec2db5d8",
  1371 => x"08802e89",
  1372 => x"38bcc408",
  1373 => x"8807bcc4",
  1374 => x"0c81fd51",
  1375 => x"a4ec2d81",
  1376 => x"fa51a4ec",
  1377 => x"2dafc304",
  1378 => x"81f551a4",
  1379 => x"ec2db5d8",
  1380 => x"08812a70",
  1381 => x"81065152",
  1382 => x"71802eaf",
  1383 => x"38bcd008",
  1384 => x"5271802e",
  1385 => x"8938ff12",
  1386 => x"bcd00cab",
  1387 => x"cb04bccc",
  1388 => x"0810bccc",
  1389 => x"08057084",
  1390 => x"29165152",
  1391 => x"88120880",
  1392 => x"2e8938ff",
  1393 => x"51881208",
  1394 => x"52712d81",
  1395 => x"f251a4ec",
  1396 => x"2db5d808",
  1397 => x"812a7081",
  1398 => x"06515271",
  1399 => x"802eb138",
  1400 => x"bccc08ff",
  1401 => x"11bcd008",
  1402 => x"56535373",
  1403 => x"72258938",
  1404 => x"8114bcd0",
  1405 => x"0cac9004",
  1406 => x"72101370",
  1407 => x"84291651",
  1408 => x"52881208",
  1409 => x"802e8938",
  1410 => x"fe518812",
  1411 => x"0852712d",
  1412 => x"81fd51a4",
  1413 => x"ec2db5d8",
  1414 => x"08812a70",
  1415 => x"81065152",
  1416 => x"71802e86",
  1417 => x"38800bbc",
  1418 => x"d00c81fa",
  1419 => x"51a4ec2d",
  1420 => x"b5d80881",
  1421 => x"2a708106",
  1422 => x"51527180",
  1423 => x"2e8938bc",
  1424 => x"cc08ff05",
  1425 => x"bcd00cbc",
  1426 => x"d0087053",
  1427 => x"5473802e",
  1428 => x"8a388c15",
  1429 => x"ff155555",
  1430 => x"accd0482",
  1431 => x"0bb5ec0c",
  1432 => x"718f06b5",
  1433 => x"e80c81eb",
  1434 => x"51a4ec2d",
  1435 => x"b5d80881",
  1436 => x"2a708106",
  1437 => x"51527180",
  1438 => x"2ead3874",
  1439 => x"08852e09",
  1440 => x"8106a438",
  1441 => x"881580f5",
  1442 => x"2dff0552",
  1443 => x"71881681",
  1444 => x"b72d7198",
  1445 => x"2b527180",
  1446 => x"25883880",
  1447 => x"0b881681",
  1448 => x"b72d7451",
  1449 => x"a5e22d81",
  1450 => x"f451a4ec",
  1451 => x"2db5d808",
  1452 => x"812a7081",
  1453 => x"06515271",
  1454 => x"802eb338",
  1455 => x"7408852e",
  1456 => x"098106aa",
  1457 => x"38881580",
  1458 => x"f52d8105",
  1459 => x"52718816",
  1460 => x"81b72d71",
  1461 => x"81ff068b",
  1462 => x"1680f52d",
  1463 => x"54527272",
  1464 => x"27873872",
  1465 => x"881681b7",
  1466 => x"2d7451a5",
  1467 => x"e22d80da",
  1468 => x"51a4ec2d",
  1469 => x"b5d80881",
  1470 => x"2a708106",
  1471 => x"51527180",
  1472 => x"2e80ff38",
  1473 => x"bcc808bc",
  1474 => x"d0085553",
  1475 => x"73802e8a",
  1476 => x"388c13ff",
  1477 => x"155553ae",
  1478 => x"8c047208",
  1479 => x"5271822e",
  1480 => x"a6387182",
  1481 => x"26893871",
  1482 => x"812ea938",
  1483 => x"af820471",
  1484 => x"832eb138",
  1485 => x"71842e09",
  1486 => x"810680c6",
  1487 => x"38881308",
  1488 => x"51a7ad2d",
  1489 => x"af8204bc",
  1490 => x"d0085188",
  1491 => x"13085271",
  1492 => x"2daf8204",
  1493 => x"810b8814",
  1494 => x"082bbcbc",
  1495 => x"0832bcbc",
  1496 => x"0caeff04",
  1497 => x"881380f5",
  1498 => x"2d81058b",
  1499 => x"1480f52d",
  1500 => x"53547174",
  1501 => x"24833880",
  1502 => x"54738814",
  1503 => x"81b72da6",
  1504 => x"922d8054",
  1505 => x"800bb5ec",
  1506 => x"0c738f06",
  1507 => x"b5e80ca0",
  1508 => x"5273bcd0",
  1509 => x"082e0981",
  1510 => x"069838bc",
  1511 => x"cc08ff05",
  1512 => x"74327009",
  1513 => x"81057072",
  1514 => x"079f2a91",
  1515 => x"71315151",
  1516 => x"53537151",
  1517 => x"82ee2d81",
  1518 => x"14548e74",
  1519 => x"25c638b5",
  1520 => x"d4085271",
  1521 => x"b5d80c02",
  1522 => x"94050d04",
  1523 => x"00ffffff",
  1524 => x"ff00ffff",
  1525 => x"ffff00ff",
  1526 => x"ffffff00",
  1527 => x"52657365",
  1528 => x"74000000",
  1529 => x"53617665",
  1530 => x"20736574",
  1531 => x"74696e67",
  1532 => x"73000000",
  1533 => x"5363616e",
  1534 => x"6c696e65",
  1535 => x"73000000",
  1536 => x"4c6f6164",
  1537 => x"20524f4d",
  1538 => x"20100000",
  1539 => x"45786974",
  1540 => x"00000000",
  1541 => x"50432045",
  1542 => x"6e67696e",
  1543 => x"65206d6f",
  1544 => x"64650000",
  1545 => x"54757262",
  1546 => x"6f677261",
  1547 => x"66782031",
  1548 => x"36206d6f",
  1549 => x"64650000",
  1550 => x"56474120",
  1551 => x"2d203331",
  1552 => x"4b487a2c",
  1553 => x"20363048",
  1554 => x"7a000000",
  1555 => x"5456202d",
  1556 => x"20343830",
  1557 => x"692c2036",
  1558 => x"30487a00",
  1559 => x"4261636b",
  1560 => x"00000000",
  1561 => x"46504741",
  1562 => x"50434520",
  1563 => x"43464700",
  1564 => x"52656164",
  1565 => x"20666169",
  1566 => x"6c65640a",
  1567 => x"00000000",
  1568 => x"4661696c",
  1569 => x"65640a00",
  1570 => x"4c6f6164",
  1571 => x"696e6720",
  1572 => x"00000000",
  1573 => x"496e6974",
  1574 => x"69616c69",
  1575 => x"7a696e67",
  1576 => x"20534420",
  1577 => x"63617264",
  1578 => x"0a000000",
  1579 => x"424f4f54",
  1580 => x"20202020",
  1581 => x"50434500",
  1582 => x"43617264",
  1583 => x"20696e69",
  1584 => x"74206661",
  1585 => x"696c6564",
  1586 => x"0a000000",
  1587 => x"4d425220",
  1588 => x"6661696c",
  1589 => x"0a000000",
  1590 => x"46415431",
  1591 => x"36202020",
  1592 => x"00000000",
  1593 => x"46415433",
  1594 => x"32202020",
  1595 => x"00000000",
  1596 => x"4e6f2070",
  1597 => x"61727469",
  1598 => x"74696f6e",
  1599 => x"20736967",
  1600 => x"0a000000",
  1601 => x"42616420",
  1602 => x"70617274",
  1603 => x"0a000000",
  1604 => x"53444843",
  1605 => x"20657272",
  1606 => x"6f72210a",
  1607 => x"00000000",
  1608 => x"53442069",
  1609 => x"6e69742e",
  1610 => x"2e2e0a00",
  1611 => x"53442063",
  1612 => x"61726420",
  1613 => x"72657365",
  1614 => x"74206661",
  1615 => x"696c6564",
  1616 => x"210a0000",
  1617 => x"57726974",
  1618 => x"65206661",
  1619 => x"696c6564",
  1620 => x"0a000000",
  1621 => x"16200000",
  1622 => x"14200000",
  1623 => x"15200000",
  1624 => x"00000002",
  1625 => x"00000002",
  1626 => x"000017dc",
  1627 => x"000004eb",
  1628 => x"00000002",
  1629 => x"000017e4",
  1630 => x"000003b3",
  1631 => x"00000003",
  1632 => x"000019cc",
  1633 => x"00000002",
  1634 => x"00000001",
  1635 => x"000017f4",
  1636 => x"00000002",
  1637 => x"00000003",
  1638 => x"000019c4",
  1639 => x"00000002",
  1640 => x"00000002",
  1641 => x"00001800",
  1642 => x"0000064b",
  1643 => x"00000002",
  1644 => x"0000180c",
  1645 => x"000012cf",
  1646 => x"00000000",
  1647 => x"00000000",
  1648 => x"00000000",
  1649 => x"00001814",
  1650 => x"00001824",
  1651 => x"00001838",
  1652 => x"0000184c",
  1653 => x"00000002",
  1654 => x"00001b0c",
  1655 => x"00000500",
  1656 => x"00000002",
  1657 => x"00001b1c",
  1658 => x"00000500",
  1659 => x"00000002",
  1660 => x"00001b2c",
  1661 => x"00000500",
  1662 => x"00000002",
  1663 => x"00001b3c",
  1664 => x"00000500",
  1665 => x"00000002",
  1666 => x"00001b4c",
  1667 => x"00000500",
  1668 => x"00000002",
  1669 => x"00001b5c",
  1670 => x"00000500",
  1671 => x"00000002",
  1672 => x"00001b6c",
  1673 => x"00000500",
  1674 => x"00000002",
  1675 => x"00001b7c",
  1676 => x"00000500",
  1677 => x"00000002",
  1678 => x"00001b8c",
  1679 => x"00000500",
  1680 => x"00000002",
  1681 => x"00001b9c",
  1682 => x"00000500",
  1683 => x"00000002",
  1684 => x"00001bac",
  1685 => x"00000500",
  1686 => x"00000002",
  1687 => x"00001bbc",
  1688 => x"00000500",
  1689 => x"00000002",
  1690 => x"00001bcc",
  1691 => x"00000500",
  1692 => x"00000004",
  1693 => x"0000185c",
  1694 => x"00001964",
  1695 => x"00000000",
  1696 => x"00000000",
  1697 => x"000005df",
  1698 => x"00000000",
  1699 => x"00000000",
  1700 => x"00000000",
  1701 => x"00000000",
  1702 => x"00000000",
  1703 => x"00000000",
  1704 => x"00000000",
  1705 => x"00000000",
  1706 => x"00000000",
  1707 => x"00000000",
  1708 => x"00000000",
  1709 => x"00000000",
  1710 => x"00000000",
  1711 => x"00000000",
  1712 => x"00000000",
  1713 => x"00000000",
  1714 => x"00000000",
  1715 => x"00000000",
  1716 => x"00000000",
  1717 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

