-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb5",
     9 => x"ac080b0b",
    10 => x"0bb5b008",
    11 => x"0b0b0bb5",
    12 => x"b4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b5b40c0b",
    16 => x"0b0bb5b0",
    17 => x"0c0b0b0b",
    18 => x"b5ac0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bafa0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b5ac70bc",
    57 => x"a0278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8cc50402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b5bc0c9f",
    65 => x"0bb5c00c",
    66 => x"a0717081",
    67 => x"055334b5",
    68 => x"c008ff05",
    69 => x"b5c00cb5",
    70 => x"c0088025",
    71 => x"eb38b5bc",
    72 => x"08ff05b5",
    73 => x"bc0cb5bc",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb5bc",
    94 => x"08258f38",
    95 => x"82b22db5",
    96 => x"bc08ff05",
    97 => x"b5bc0c82",
    98 => x"f404b5bc",
    99 => x"08b5c008",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b5bc08",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b5",
   108 => x"c0088105",
   109 => x"b5c00cb5",
   110 => x"c008519f",
   111 => x"7125e238",
   112 => x"800bb5c0",
   113 => x"0cb5bc08",
   114 => x"8105b5bc",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b5c00881",
   120 => x"05b5c00c",
   121 => x"b5c008a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b5c00cb5",
   125 => x"bc088105",
   126 => x"b5bc0c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb5",
   155 => x"c40cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb5c4",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b5c40884",
   167 => x"07b5c40c",
   168 => x"5573842b",
   169 => x"87e87125",
   170 => x"83713170",
   171 => x"0b0b0bb2",
   172 => x"b40c8171",
   173 => x"2bf6880c",
   174 => x"fea413ff",
   175 => x"122c7888",
   176 => x"29ff9405",
   177 => x"70812cb5",
   178 => x"c4085258",
   179 => x"52555152",
   180 => x"5476802e",
   181 => x"85387081",
   182 => x"075170f6",
   183 => x"940c7109",
   184 => x"8105f680",
   185 => x"0c720981",
   186 => x"05f6840c",
   187 => x"0294050d",
   188 => x"0402f405",
   189 => x"0d745372",
   190 => x"70810554",
   191 => x"80f52d52",
   192 => x"71802e89",
   193 => x"38715182",
   194 => x"ee2d85f7",
   195 => x"04028c05",
   196 => x"0d0402f4",
   197 => x"050d7470",
   198 => x"8206bc88",
   199 => x"0cb2d071",
   200 => x"81065454",
   201 => x"51718814",
   202 => x"81b72d70",
   203 => x"822a7081",
   204 => x"06515170",
   205 => x"941481b7",
   206 => x"2d70b5ac",
   207 => x"0c028c05",
   208 => x"0d0402f4",
   209 => x"050db0b8",
   210 => x"52b5cc51",
   211 => x"95de2db5",
   212 => x"ac08802e",
   213 => x"9538b7a8",
   214 => x"52b5cc51",
   215 => x"98942db7",
   216 => x"a80870fe",
   217 => x"c00c5186",
   218 => x"922d028c",
   219 => x"050d0402",
   220 => x"f8050dbc",
   221 => x"88088206",
   222 => x"b2d80b80",
   223 => x"f52d5252",
   224 => x"70802e85",
   225 => x"38718107",
   226 => x"52b2f00b",
   227 => x"80f52d51",
   228 => x"70802e85",
   229 => x"38718407",
   230 => x"5271b5ac",
   231 => x"0c028805",
   232 => x"0d0402f0",
   233 => x"050d86ef",
   234 => x"2db5ac08",
   235 => x"b0b853b5",
   236 => x"cc525395",
   237 => x"de2db5ac",
   238 => x"08802ea3",
   239 => x"3872b7a8",
   240 => x"0cb7ac54",
   241 => x"80fd5380",
   242 => x"74708405",
   243 => x"560cff13",
   244 => x"53728025",
   245 => x"f238b7a8",
   246 => x"52b5cc51",
   247 => x"98ba2d02",
   248 => x"90050d04",
   249 => x"02d8050d",
   250 => x"810bfec4",
   251 => x"0c840bfe",
   252 => x"c40c7b52",
   253 => x"b5cc5195",
   254 => x"de2db5ac",
   255 => x"0853b5ac",
   256 => x"08802e81",
   257 => x"ba38b5d0",
   258 => x"0856800b",
   259 => x"ff175859",
   260 => x"76792e8b",
   261 => x"38811977",
   262 => x"812a5859",
   263 => x"76f738f7",
   264 => x"19769fff",
   265 => x"06545972",
   266 => x"802e8b38",
   267 => x"fc8016b5",
   268 => x"cc525697",
   269 => x"e72d8076",
   270 => x"2580fa38",
   271 => x"78527651",
   272 => x"84802db7",
   273 => x"a852b5cc",
   274 => x"5198942d",
   275 => x"b5ac0853",
   276 => x"b5ac0880",
   277 => x"2e80c838",
   278 => x"b7a85a80",
   279 => x"58898c04",
   280 => x"79708405",
   281 => x"5b087083",
   282 => x"fe800671",
   283 => x"882b83fe",
   284 => x"80067188",
   285 => x"2a077288",
   286 => x"2a83fe80",
   287 => x"0673982a",
   288 => x"07fec80c",
   289 => x"fec80c56",
   290 => x"84195953",
   291 => x"75538480",
   292 => x"76258438",
   293 => x"84805372",
   294 => x"7824c538",
   295 => x"89a504b0",
   296 => x"c45189c2",
   297 => x"04b5cc51",
   298 => x"97e72dfc",
   299 => x"80168118",
   300 => x"585688b6",
   301 => x"04820bfe",
   302 => x"c40c8153",
   303 => x"89c504b0",
   304 => x"d45185f1",
   305 => x"2d72b5ac",
   306 => x"0c02a805",
   307 => x"0d0402fc",
   308 => x"050da5a3",
   309 => x"2dfec451",
   310 => x"81710c82",
   311 => x"710c0284",
   312 => x"050d0402",
   313 => x"f4050d74",
   314 => x"10157084",
   315 => x"29b3ac05",
   316 => x"70085551",
   317 => x"5272802e",
   318 => x"9b387280",
   319 => x"f52d5271",
   320 => x"802e9138",
   321 => x"b0dc5185",
   322 => x"f12d7251",
   323 => x"85f12d72",
   324 => x"5187e42d",
   325 => x"b2b851a7",
   326 => x"812da5a3",
   327 => x"2d805184",
   328 => x"e52d028c",
   329 => x"050d0402",
   330 => x"e8050d80",
   331 => x"70565675",
   332 => x"b4dc0825",
   333 => x"af38bbb4",
   334 => x"08762ea8",
   335 => x"38745195",
   336 => x"892db5ac",
   337 => x"08098105",
   338 => x"70b5ac08",
   339 => x"079f2a77",
   340 => x"05811757",
   341 => x"575275b4",
   342 => x"dc082588",
   343 => x"38bbb408",
   344 => x"7526da38",
   345 => x"805674bb",
   346 => x"b4082780",
   347 => x"d0387451",
   348 => x"95892d75",
   349 => x"842b52b5",
   350 => x"ac08802e",
   351 => x"ae38b5d8",
   352 => x"128117b5",
   353 => x"ac085657",
   354 => x"528a5373",
   355 => x"70810555",
   356 => x"80f52d72",
   357 => x"70810554",
   358 => x"81b72dff",
   359 => x"13537280",
   360 => x"25e93880",
   361 => x"7281b72d",
   362 => x"8bb404b5",
   363 => x"ac08b5d8",
   364 => x"1381b72d",
   365 => x"8115558b",
   366 => x"7625ffaa",
   367 => x"38029805",
   368 => x"0d0402fc",
   369 => x"050d7251",
   370 => x"70fd2ead",
   371 => x"3870fd24",
   372 => x"8a3870fc",
   373 => x"2e80c438",
   374 => x"8ca30470",
   375 => x"fe2eb138",
   376 => x"70ff2e09",
   377 => x"8106bc38",
   378 => x"b4dc0851",
   379 => x"70802eb3",
   380 => x"38ff11b4",
   381 => x"dc0c8ca3",
   382 => x"04b4dc08",
   383 => x"f00570b4",
   384 => x"dc0c5170",
   385 => x"80259c38",
   386 => x"800bb4dc",
   387 => x"0c8ca304",
   388 => x"b4dc0881",
   389 => x"05b4dc0c",
   390 => x"8ca304b4",
   391 => x"dc089005",
   392 => x"b4dc0c8a",
   393 => x"a72da5e6",
   394 => x"2d028405",
   395 => x"0d0402fc",
   396 => x"050d800b",
   397 => x"b4dc0c8a",
   398 => x"a72db3a8",
   399 => x"51a7812d",
   400 => x"0284050d",
   401 => x"0402f405",
   402 => x"0d805186",
   403 => x"922d810b",
   404 => x"fec40c80",
   405 => x"0bfec00c",
   406 => x"840bfec4",
   407 => x"0c830bfe",
   408 => x"cc0ca2f1",
   409 => x"2da5842d",
   410 => x"a2d62da2",
   411 => x"d62d81f7",
   412 => x"2d815184",
   413 => x"e52da2d6",
   414 => x"2da2d62d",
   415 => x"815184e5",
   416 => x"2db0e851",
   417 => x"85f12d84",
   418 => x"529ced2d",
   419 => x"8ef72db5",
   420 => x"ac08802e",
   421 => x"8638fe52",
   422 => x"8da304ff",
   423 => x"12527180",
   424 => x"24e73871",
   425 => x"802e8181",
   426 => x"3886c22d",
   427 => x"b1805187",
   428 => x"e42db5ac",
   429 => x"08802e8f",
   430 => x"38b2b851",
   431 => x"a7812d80",
   432 => x"5184e52d",
   433 => x"8dd104b5",
   434 => x"ac08518c",
   435 => x"ae2da590",
   436 => x"2da3892d",
   437 => x"a7912db5",
   438 => x"ac08bc8c",
   439 => x"08882bbc",
   440 => x"900807fe",
   441 => x"d80c5386",
   442 => x"ef2db5ac",
   443 => x"08b5c808",
   444 => x"2ea238b5",
   445 => x"ac08b5c8",
   446 => x"0cb5ac08",
   447 => x"fec00c84",
   448 => x"52725184",
   449 => x"e52da2d6",
   450 => x"2da2d62d",
   451 => x"ff125271",
   452 => x"8025ee38",
   453 => x"72802e89",
   454 => x"388a0bfe",
   455 => x"c40c8dd1",
   456 => x"04820bfe",
   457 => x"c40c8dd1",
   458 => x"04b18c51",
   459 => x"85f12d80",
   460 => x"0bb5ac0c",
   461 => x"028c050d",
   462 => x"0402e805",
   463 => x"0d77797b",
   464 => x"58555580",
   465 => x"53727625",
   466 => x"a3387470",
   467 => x"81055680",
   468 => x"f52d7470",
   469 => x"81055680",
   470 => x"f52d5252",
   471 => x"71712e86",
   472 => x"3881518e",
   473 => x"ee048113",
   474 => x"538ec504",
   475 => x"805170b5",
   476 => x"ac0c0298",
   477 => x"050d0402",
   478 => x"d8050d80",
   479 => x"0bbbb00c",
   480 => x"b7a85280",
   481 => x"519fd52d",
   482 => x"b5ac0854",
   483 => x"b5ac088c",
   484 => x"38b1a051",
   485 => x"85f12d73",
   486 => x"55949204",
   487 => x"8056810b",
   488 => x"bbd40c88",
   489 => x"53b1ac52",
   490 => x"b7de518e",
   491 => x"b92db5ac",
   492 => x"08762e09",
   493 => x"81068738",
   494 => x"b5ac08bb",
   495 => x"d40c8853",
   496 => x"b1b852b7",
   497 => x"fa518eb9",
   498 => x"2db5ac08",
   499 => x"8738b5ac",
   500 => x"08bbd40c",
   501 => x"bbd40880",
   502 => x"2e80f638",
   503 => x"baee0b80",
   504 => x"f52dbaef",
   505 => x"0b80f52d",
   506 => x"71982b71",
   507 => x"902b07ba",
   508 => x"f00b80f5",
   509 => x"2d70882b",
   510 => x"7207baf1",
   511 => x"0b80f52d",
   512 => x"7107bba6",
   513 => x"0b80f52d",
   514 => x"bba70b80",
   515 => x"f52d7188",
   516 => x"2b07535f",
   517 => x"54525a56",
   518 => x"57557381",
   519 => x"abaa2e09",
   520 => x"81068d38",
   521 => x"7551a0f0",
   522 => x"2db5ac08",
   523 => x"5690bd04",
   524 => x"7382d4d5",
   525 => x"2e8738b1",
   526 => x"c45190fe",
   527 => x"04b7a852",
   528 => x"75519fd5",
   529 => x"2db5ac08",
   530 => x"55b5ac08",
   531 => x"802e83c2",
   532 => x"388853b1",
   533 => x"b852b7fa",
   534 => x"518eb92d",
   535 => x"b5ac0889",
   536 => x"38810bbb",
   537 => x"b00c9184",
   538 => x"048853b1",
   539 => x"ac52b7de",
   540 => x"518eb92d",
   541 => x"b5ac0880",
   542 => x"2e8a38b1",
   543 => x"d85185f1",
   544 => x"2d91de04",
   545 => x"bba60b80",
   546 => x"f52d5473",
   547 => x"80d52e09",
   548 => x"810680ca",
   549 => x"38bba70b",
   550 => x"80f52d54",
   551 => x"7381aa2e",
   552 => x"098106ba",
   553 => x"38800bb7",
   554 => x"a80b80f5",
   555 => x"2d565474",
   556 => x"81e92e83",
   557 => x"38815474",
   558 => x"81eb2e8c",
   559 => x"38805573",
   560 => x"752e0981",
   561 => x"0682cb38",
   562 => x"b7b30b80",
   563 => x"f52d5574",
   564 => x"8d38b7b4",
   565 => x"0b80f52d",
   566 => x"5473822e",
   567 => x"86388055",
   568 => x"949204b7",
   569 => x"b50b80f5",
   570 => x"2d70bba8",
   571 => x"0cff05bb",
   572 => x"ac0cb7b6",
   573 => x"0b80f52d",
   574 => x"b7b70b80",
   575 => x"f52d5876",
   576 => x"05778280",
   577 => x"290570bb",
   578 => x"b80cb7b8",
   579 => x"0b80f52d",
   580 => x"70bbcc0c",
   581 => x"bbb00859",
   582 => x"57587680",
   583 => x"2e81a338",
   584 => x"8853b1b8",
   585 => x"52b7fa51",
   586 => x"8eb92db5",
   587 => x"ac0881e2",
   588 => x"38bba808",
   589 => x"70842bbb",
   590 => x"b40c70bb",
   591 => x"c80cb7cd",
   592 => x"0b80f52d",
   593 => x"b7cc0b80",
   594 => x"f52d7182",
   595 => x"802905b7",
   596 => x"ce0b80f5",
   597 => x"2d708480",
   598 => x"802912b7",
   599 => x"cf0b80f5",
   600 => x"2d708180",
   601 => x"0a291270",
   602 => x"bbd00cbb",
   603 => x"cc087129",
   604 => x"bbb80805",
   605 => x"70bbbc0c",
   606 => x"b7d50b80",
   607 => x"f52db7d4",
   608 => x"0b80f52d",
   609 => x"71828029",
   610 => x"05b7d60b",
   611 => x"80f52d70",
   612 => x"84808029",
   613 => x"12b7d70b",
   614 => x"80f52d70",
   615 => x"982b81f0",
   616 => x"0a067205",
   617 => x"70bbc00c",
   618 => x"fe117e29",
   619 => x"7705bbc4",
   620 => x"0c525952",
   621 => x"43545e51",
   622 => x"5259525d",
   623 => x"57595794",
   624 => x"9004b7ba",
   625 => x"0b80f52d",
   626 => x"b7b90b80",
   627 => x"f52d7182",
   628 => x"80290570",
   629 => x"bbb40c70",
   630 => x"a02983ff",
   631 => x"0570892a",
   632 => x"70bbc80c",
   633 => x"b7bf0b80",
   634 => x"f52db7be",
   635 => x"0b80f52d",
   636 => x"71828029",
   637 => x"0570bbd0",
   638 => x"0c7b7129",
   639 => x"1e70bbc4",
   640 => x"0c7dbbc0",
   641 => x"0c7305bb",
   642 => x"bc0c555e",
   643 => x"51515555",
   644 => x"815574b5",
   645 => x"ac0c02a8",
   646 => x"050d0402",
   647 => x"ec050d76",
   648 => x"70872c71",
   649 => x"80ff0655",
   650 => x"5654bbb0",
   651 => x"088a3873",
   652 => x"882c7481",
   653 => x"ff065455",
   654 => x"b7a852bb",
   655 => x"b8081551",
   656 => x"9fd52db5",
   657 => x"ac0854b5",
   658 => x"ac08802e",
   659 => x"b338bbb0",
   660 => x"08802e98",
   661 => x"38728429",
   662 => x"b7a80570",
   663 => x"085253a0",
   664 => x"f02db5ac",
   665 => x"08f00a06",
   666 => x"5394fe04",
   667 => x"7210b7a8",
   668 => x"057080e0",
   669 => x"2d5253a1",
   670 => x"a02db5ac",
   671 => x"08537254",
   672 => x"73b5ac0c",
   673 => x"0294050d",
   674 => x"0402ec05",
   675 => x"0d767084",
   676 => x"2cbbc408",
   677 => x"05718f06",
   678 => x"52555372",
   679 => x"8938b7a8",
   680 => x"5273519f",
   681 => x"d52d72a0",
   682 => x"29b7a805",
   683 => x"54807480",
   684 => x"f52d5455",
   685 => x"72752e83",
   686 => x"38815572",
   687 => x"81e52e93",
   688 => x"3874802e",
   689 => x"8e388b14",
   690 => x"80f52d98",
   691 => x"06537280",
   692 => x"2e833880",
   693 => x"5473b5ac",
   694 => x"0c029405",
   695 => x"0d0402cc",
   696 => x"050d7e60",
   697 => x"5e5a800b",
   698 => x"bbc008bb",
   699 => x"c408595c",
   700 => x"568058bb",
   701 => x"b408782e",
   702 => x"81ae3877",
   703 => x"8f06a017",
   704 => x"5754738f",
   705 => x"38b7a852",
   706 => x"76518117",
   707 => x"579fd52d",
   708 => x"b7a85680",
   709 => x"7680f52d",
   710 => x"56547474",
   711 => x"2e833881",
   712 => x"547481e5",
   713 => x"2e80f638",
   714 => x"81707506",
   715 => x"555c7380",
   716 => x"2e80ea38",
   717 => x"8b1680f5",
   718 => x"2d980659",
   719 => x"7880de38",
   720 => x"8b537c52",
   721 => x"75518eb9",
   722 => x"2db5ac08",
   723 => x"80cf389c",
   724 => x"160851a0",
   725 => x"f02db5ac",
   726 => x"08841b0c",
   727 => x"9a1680e0",
   728 => x"2d51a1a0",
   729 => x"2db5ac08",
   730 => x"b5ac0888",
   731 => x"1c0cb5ac",
   732 => x"085555bb",
   733 => x"b008802e",
   734 => x"98389416",
   735 => x"80e02d51",
   736 => x"a1a02db5",
   737 => x"ac08902b",
   738 => x"83fff00a",
   739 => x"06701651",
   740 => x"5473881b",
   741 => x"0c787a0c",
   742 => x"7b5497de",
   743 => x"04811858",
   744 => x"bbb40878",
   745 => x"26fed438",
   746 => x"bbb00880",
   747 => x"2eae387a",
   748 => x"51949b2d",
   749 => x"b5ac08b5",
   750 => x"ac0880ff",
   751 => x"fffff806",
   752 => x"555b7380",
   753 => x"fffffff8",
   754 => x"2e9238b5",
   755 => x"ac08fe05",
   756 => x"bba80829",
   757 => x"bbbc0805",
   758 => x"5795f104",
   759 => x"805473b5",
   760 => x"ac0c02b4",
   761 => x"050d0402",
   762 => x"f4050d74",
   763 => x"70088105",
   764 => x"710c7008",
   765 => x"bbac0806",
   766 => x"5353718e",
   767 => x"38881308",
   768 => x"51949b2d",
   769 => x"b5ac0888",
   770 => x"140c810b",
   771 => x"b5ac0c02",
   772 => x"8c050d04",
   773 => x"02f0050d",
   774 => x"75881108",
   775 => x"fe05bba8",
   776 => x"0829bbbc",
   777 => x"08117208",
   778 => x"bbac0806",
   779 => x"05795553",
   780 => x"54549fd5",
   781 => x"2d029005",
   782 => x"0d0402f0",
   783 => x"050d7588",
   784 => x"1108fe05",
   785 => x"bba80829",
   786 => x"bbbc0811",
   787 => x"7208bbac",
   788 => x"08060579",
   789 => x"55535454",
   790 => x"9e952d02",
   791 => x"90050d04",
   792 => x"02f4050d",
   793 => x"d45281ff",
   794 => x"720c7108",
   795 => x"5381ff72",
   796 => x"0c72882b",
   797 => x"83fe8006",
   798 => x"72087081",
   799 => x"ff065152",
   800 => x"5381ff72",
   801 => x"0c727107",
   802 => x"882b7208",
   803 => x"7081ff06",
   804 => x"51525381",
   805 => x"ff720c72",
   806 => x"7107882b",
   807 => x"72087081",
   808 => x"ff067207",
   809 => x"b5ac0c52",
   810 => x"53028c05",
   811 => x"0d0402f4",
   812 => x"050d7476",
   813 => x"7181ff06",
   814 => x"d40c5353",
   815 => x"bbd80885",
   816 => x"3871892b",
   817 => x"5271982a",
   818 => x"d40c7190",
   819 => x"2a7081ff",
   820 => x"06d40c51",
   821 => x"71882a70",
   822 => x"81ff06d4",
   823 => x"0c517181",
   824 => x"ff06d40c",
   825 => x"72902a70",
   826 => x"81ff06d4",
   827 => x"0c51d408",
   828 => x"7081ff06",
   829 => x"515182b8",
   830 => x"bf527081",
   831 => x"ff2e0981",
   832 => x"06943881",
   833 => x"ff0bd40c",
   834 => x"d4087081",
   835 => x"ff06ff14",
   836 => x"54515171",
   837 => x"e53870b5",
   838 => x"ac0c028c",
   839 => x"050d0402",
   840 => x"fc050d81",
   841 => x"c75181ff",
   842 => x"0bd40cff",
   843 => x"11517080",
   844 => x"25f43802",
   845 => x"84050d04",
   846 => x"02f0050d",
   847 => x"9a9f2d8f",
   848 => x"cf538052",
   849 => x"87fc80f7",
   850 => x"5199ae2d",
   851 => x"b5ac0854",
   852 => x"b5ac0881",
   853 => x"2e098106",
   854 => x"a33881ff",
   855 => x"0bd40c82",
   856 => x"0a52849c",
   857 => x"80e95199",
   858 => x"ae2db5ac",
   859 => x"088b3881",
   860 => x"ff0bd40c",
   861 => x"73539b82",
   862 => x"049a9f2d",
   863 => x"ff135372",
   864 => x"c13872b5",
   865 => x"ac0c0290",
   866 => x"050d0402",
   867 => x"f4050d81",
   868 => x"ff0bd40c",
   869 => x"93538052",
   870 => x"87fc80c1",
   871 => x"5199ae2d",
   872 => x"b5ac088b",
   873 => x"3881ff0b",
   874 => x"d40c8153",
   875 => x"9bb8049a",
   876 => x"9f2dff13",
   877 => x"5372df38",
   878 => x"72b5ac0c",
   879 => x"028c050d",
   880 => x"0402f005",
   881 => x"0d9a9f2d",
   882 => x"83aa5284",
   883 => x"9c80c851",
   884 => x"99ae2db5",
   885 => x"ac08812e",
   886 => x"09810692",
   887 => x"3898e02d",
   888 => x"b5ac0883",
   889 => x"ffff0653",
   890 => x"7283aa2e",
   891 => x"97389b8b",
   892 => x"2d9bff04",
   893 => x"81549ce4",
   894 => x"04b1e451",
   895 => x"85f12d80",
   896 => x"549ce404",
   897 => x"81ff0bd4",
   898 => x"0cb1539a",
   899 => x"b82db5ac",
   900 => x"08802e80",
   901 => x"c0388052",
   902 => x"87fc80fa",
   903 => x"5199ae2d",
   904 => x"b5ac08b1",
   905 => x"3881ff0b",
   906 => x"d40cd408",
   907 => x"5381ff0b",
   908 => x"d40c81ff",
   909 => x"0bd40c81",
   910 => x"ff0bd40c",
   911 => x"81ff0bd4",
   912 => x"0c72862a",
   913 => x"708106b5",
   914 => x"ac085651",
   915 => x"5372802e",
   916 => x"93389bf4",
   917 => x"0472822e",
   918 => x"ff9f38ff",
   919 => x"135372ff",
   920 => x"aa387254",
   921 => x"73b5ac0c",
   922 => x"0290050d",
   923 => x"0402f005",
   924 => x"0d810bbb",
   925 => x"d80c8454",
   926 => x"d008708f",
   927 => x"2a708106",
   928 => x"51515372",
   929 => x"f33872d0",
   930 => x"0c9a9f2d",
   931 => x"b1f45185",
   932 => x"f12dd008",
   933 => x"708f2a70",
   934 => x"81065151",
   935 => x"5372f338",
   936 => x"810bd00c",
   937 => x"b1538052",
   938 => x"84d480c0",
   939 => x"5199ae2d",
   940 => x"b5ac0881",
   941 => x"2ea13872",
   942 => x"822e0981",
   943 => x"068c38b2",
   944 => x"805185f1",
   945 => x"2d80539e",
   946 => x"8c04ff13",
   947 => x"5372d738",
   948 => x"ff145473",
   949 => x"ffa2389b",
   950 => x"c12db5ac",
   951 => x"08bbd80c",
   952 => x"b5ac088b",
   953 => x"38815287",
   954 => x"fc80d051",
   955 => x"99ae2d81",
   956 => x"ff0bd40c",
   957 => x"d008708f",
   958 => x"2a708106",
   959 => x"51515372",
   960 => x"f33872d0",
   961 => x"0c81ff0b",
   962 => x"d40c8153",
   963 => x"72b5ac0c",
   964 => x"0290050d",
   965 => x"0402e805",
   966 => x"0d785681",
   967 => x"ff0bd40c",
   968 => x"d008708f",
   969 => x"2a708106",
   970 => x"51515372",
   971 => x"f3388281",
   972 => x"0bd00c81",
   973 => x"ff0bd40c",
   974 => x"775287fc",
   975 => x"80d85199",
   976 => x"ae2db5ac",
   977 => x"08802e8c",
   978 => x"38b29851",
   979 => x"85f12d81",
   980 => x"539fcc04",
   981 => x"81ff0bd4",
   982 => x"0c81fe0b",
   983 => x"d40c80ff",
   984 => x"55757084",
   985 => x"05570870",
   986 => x"982ad40c",
   987 => x"70902c70",
   988 => x"81ff06d4",
   989 => x"0c547088",
   990 => x"2c7081ff",
   991 => x"06d40c54",
   992 => x"7081ff06",
   993 => x"d40c54ff",
   994 => x"15557480",
   995 => x"25d33881",
   996 => x"ff0bd40c",
   997 => x"81ff0bd4",
   998 => x"0c81ff0b",
   999 => x"d40c868d",
  1000 => x"a05481ff",
  1001 => x"0bd40cd4",
  1002 => x"0881ff06",
  1003 => x"55748738",
  1004 => x"ff145473",
  1005 => x"ed3881ff",
  1006 => x"0bd40cd0",
  1007 => x"08708f2a",
  1008 => x"70810651",
  1009 => x"515372f3",
  1010 => x"3872d00c",
  1011 => x"72b5ac0c",
  1012 => x"0298050d",
  1013 => x"0402e805",
  1014 => x"0d785580",
  1015 => x"5681ff0b",
  1016 => x"d40cd008",
  1017 => x"708f2a70",
  1018 => x"81065151",
  1019 => x"5372f338",
  1020 => x"82810bd0",
  1021 => x"0c81ff0b",
  1022 => x"d40c7752",
  1023 => x"87fc80d1",
  1024 => x"5199ae2d",
  1025 => x"80dbc6df",
  1026 => x"54b5ac08",
  1027 => x"802e8a38",
  1028 => x"b0c45185",
  1029 => x"f12da0e7",
  1030 => x"0481ff0b",
  1031 => x"d40cd408",
  1032 => x"7081ff06",
  1033 => x"51537281",
  1034 => x"fe2e0981",
  1035 => x"069d3880",
  1036 => x"ff5398e0",
  1037 => x"2db5ac08",
  1038 => x"75708405",
  1039 => x"570cff13",
  1040 => x"53728025",
  1041 => x"ed388156",
  1042 => x"a0d104ff",
  1043 => x"145473c9",
  1044 => x"3881ff0b",
  1045 => x"d40cd008",
  1046 => x"708f2a70",
  1047 => x"81065151",
  1048 => x"5372f338",
  1049 => x"72d00c75",
  1050 => x"b5ac0c02",
  1051 => x"98050d04",
  1052 => x"02f4050d",
  1053 => x"7470882a",
  1054 => x"83fe8006",
  1055 => x"7072982a",
  1056 => x"0772882b",
  1057 => x"87fc8080",
  1058 => x"0673982b",
  1059 => x"81f00a06",
  1060 => x"71730707",
  1061 => x"b5ac0c56",
  1062 => x"51535102",
  1063 => x"8c050d04",
  1064 => x"02f8050d",
  1065 => x"028e0580",
  1066 => x"f52d7488",
  1067 => x"2b077083",
  1068 => x"ffff06b5",
  1069 => x"ac0c5102",
  1070 => x"88050d04",
  1071 => x"02fc050d",
  1072 => x"72518071",
  1073 => x"0c800b84",
  1074 => x"120c0284",
  1075 => x"050d0402",
  1076 => x"f0050d75",
  1077 => x"70088412",
  1078 => x"08535353",
  1079 => x"ff547171",
  1080 => x"2ea838a5",
  1081 => x"8a2d8413",
  1082 => x"08708429",
  1083 => x"14881170",
  1084 => x"087081ff",
  1085 => x"06841808",
  1086 => x"81118706",
  1087 => x"841a0c53",
  1088 => x"51555151",
  1089 => x"51a5842d",
  1090 => x"715473b5",
  1091 => x"ac0c0290",
  1092 => x"050d0402",
  1093 => x"f8050da5",
  1094 => x"8a2de008",
  1095 => x"708b2a70",
  1096 => x"81065152",
  1097 => x"5270802e",
  1098 => x"9d38bbdc",
  1099 => x"08708429",
  1100 => x"bbe40573",
  1101 => x"81ff0671",
  1102 => x"0c5151bb",
  1103 => x"dc088111",
  1104 => x"8706bbdc",
  1105 => x"0c51800b",
  1106 => x"bc840ca4",
  1107 => x"fd2da584",
  1108 => x"2d028805",
  1109 => x"0d0402fc",
  1110 => x"050da58a",
  1111 => x"2d810bbc",
  1112 => x"840ca584",
  1113 => x"2dbc8408",
  1114 => x"5170fa38",
  1115 => x"0284050d",
  1116 => x"0402fc05",
  1117 => x"0dbbdc51",
  1118 => x"a1bc2da2",
  1119 => x"9351a4f9",
  1120 => x"2da4a32d",
  1121 => x"0284050d",
  1122 => x"0402f405",
  1123 => x"0da48b04",
  1124 => x"b5ac0881",
  1125 => x"f02e0981",
  1126 => x"06893881",
  1127 => x"0bb5a00c",
  1128 => x"a48b04b5",
  1129 => x"ac0881e0",
  1130 => x"2e098106",
  1131 => x"8938810b",
  1132 => x"b5a40ca4",
  1133 => x"8b04b5ac",
  1134 => x"0852b5a4",
  1135 => x"08802e88",
  1136 => x"38b5ac08",
  1137 => x"81800552",
  1138 => x"71842c72",
  1139 => x"8f065353",
  1140 => x"b5a00880",
  1141 => x"2e993872",
  1142 => x"8429b4e0",
  1143 => x"05721381",
  1144 => x"712b7009",
  1145 => x"73080673",
  1146 => x"0c515353",
  1147 => x"a4810472",
  1148 => x"8429b4e0",
  1149 => x"05721383",
  1150 => x"712b7208",
  1151 => x"07720c53",
  1152 => x"53800bb5",
  1153 => x"a40c800b",
  1154 => x"b5a00cbb",
  1155 => x"dc51a1cf",
  1156 => x"2db5ac08",
  1157 => x"ff24fef8",
  1158 => x"38800bb5",
  1159 => x"ac0c028c",
  1160 => x"050d0402",
  1161 => x"f8050db4",
  1162 => x"e0528f51",
  1163 => x"80727084",
  1164 => x"05540cff",
  1165 => x"11517080",
  1166 => x"25f23802",
  1167 => x"88050d04",
  1168 => x"02f0050d",
  1169 => x"7551a58a",
  1170 => x"2d70822c",
  1171 => x"fc06b4e0",
  1172 => x"1172109e",
  1173 => x"06710870",
  1174 => x"722a7083",
  1175 => x"0682742b",
  1176 => x"70097406",
  1177 => x"760c5451",
  1178 => x"56575351",
  1179 => x"53a5842d",
  1180 => x"71b5ac0c",
  1181 => x"0290050d",
  1182 => x"0471980c",
  1183 => x"04ffb008",
  1184 => x"b5ac0c04",
  1185 => x"810bffb0",
  1186 => x"0c04800b",
  1187 => x"ffb00c04",
  1188 => x"02fc050d",
  1189 => x"810bb5a8",
  1190 => x"0c815184",
  1191 => x"e52d0284",
  1192 => x"050d0402",
  1193 => x"fc050d80",
  1194 => x"0bb5a80c",
  1195 => x"805184e5",
  1196 => x"2d028405",
  1197 => x"0d0402ec",
  1198 => x"050d7654",
  1199 => x"8052870b",
  1200 => x"881580f5",
  1201 => x"2d565374",
  1202 => x"72248338",
  1203 => x"a0537251",
  1204 => x"82ee2d81",
  1205 => x"128b1580",
  1206 => x"f52d5452",
  1207 => x"727225de",
  1208 => x"38029405",
  1209 => x"0d0402f0",
  1210 => x"050dbc94",
  1211 => x"085481f7",
  1212 => x"2d800bbc",
  1213 => x"980c7308",
  1214 => x"802e8180",
  1215 => x"38820bb5",
  1216 => x"c00cbc98",
  1217 => x"088f06b5",
  1218 => x"bc0c7308",
  1219 => x"5271832e",
  1220 => x"96387183",
  1221 => x"26893871",
  1222 => x"812eaf38",
  1223 => x"a6e70471",
  1224 => x"852e9f38",
  1225 => x"a6e70488",
  1226 => x"1480f52d",
  1227 => x"841508b2",
  1228 => x"a8535452",
  1229 => x"85f12d71",
  1230 => x"84291370",
  1231 => x"085252a6",
  1232 => x"eb047351",
  1233 => x"a5b62da6",
  1234 => x"e704bc88",
  1235 => x"08881508",
  1236 => x"2c708106",
  1237 => x"51527180",
  1238 => x"2e8738b2",
  1239 => x"ac51a6e4",
  1240 => x"04b2b051",
  1241 => x"85f12d84",
  1242 => x"14085185",
  1243 => x"f12dbc98",
  1244 => x"088105bc",
  1245 => x"980c8c14",
  1246 => x"54a5f604",
  1247 => x"0290050d",
  1248 => x"0471bc94",
  1249 => x"0ca5e62d",
  1250 => x"bc9808ff",
  1251 => x"05bc9c0c",
  1252 => x"0402ec05",
  1253 => x"0dbc9408",
  1254 => x"5580f851",
  1255 => x"a4c02db5",
  1256 => x"ac08812a",
  1257 => x"70810651",
  1258 => x"52719b38",
  1259 => x"8751a4c0",
  1260 => x"2db5ac08",
  1261 => x"812a7081",
  1262 => x"06515271",
  1263 => x"802eb138",
  1264 => x"a7c604a3",
  1265 => x"892d8751",
  1266 => x"a4c02db5",
  1267 => x"ac08f438",
  1268 => x"a7d604a3",
  1269 => x"892d80f8",
  1270 => x"51a4c02d",
  1271 => x"b5ac08f3",
  1272 => x"38b5a808",
  1273 => x"813270b5",
  1274 => x"a80c7052",
  1275 => x"5284e52d",
  1276 => x"800bbc8c",
  1277 => x"0c800bbc",
  1278 => x"900cb5a8",
  1279 => x"0882dd38",
  1280 => x"80da51a4",
  1281 => x"c02db5ac",
  1282 => x"08802e8a",
  1283 => x"38bc8c08",
  1284 => x"818007bc",
  1285 => x"8c0c80d9",
  1286 => x"51a4c02d",
  1287 => x"b5ac0880",
  1288 => x"2e8a38bc",
  1289 => x"8c0880c0",
  1290 => x"07bc8c0c",
  1291 => x"819451a4",
  1292 => x"c02db5ac",
  1293 => x"08802e89",
  1294 => x"38bc8c08",
  1295 => x"9007bc8c",
  1296 => x"0c819151",
  1297 => x"a4c02db5",
  1298 => x"ac08802e",
  1299 => x"8938bc8c",
  1300 => x"08a007bc",
  1301 => x"8c0c81f5",
  1302 => x"51a4c02d",
  1303 => x"b5ac0880",
  1304 => x"2e8938bc",
  1305 => x"8c088107",
  1306 => x"bc8c0c81",
  1307 => x"f251a4c0",
  1308 => x"2db5ac08",
  1309 => x"802e8938",
  1310 => x"bc8c0882",
  1311 => x"07bc8c0c",
  1312 => x"81eb51a4",
  1313 => x"c02db5ac",
  1314 => x"08802e89",
  1315 => x"38bc8c08",
  1316 => x"8407bc8c",
  1317 => x"0c81f451",
  1318 => x"a4c02db5",
  1319 => x"ac08802e",
  1320 => x"8938bc8c",
  1321 => x"088807bc",
  1322 => x"8c0c80d8",
  1323 => x"51a4c02d",
  1324 => x"b5ac0880",
  1325 => x"2e8a38bc",
  1326 => x"90088180",
  1327 => x"07bc900c",
  1328 => x"9251a4c0",
  1329 => x"2db5ac08",
  1330 => x"802e8a38",
  1331 => x"bc900880",
  1332 => x"c007bc90",
  1333 => x"0c9451a4",
  1334 => x"c02db5ac",
  1335 => x"08802e89",
  1336 => x"38bc9008",
  1337 => x"9007bc90",
  1338 => x"0c9151a4",
  1339 => x"c02db5ac",
  1340 => x"08802e89",
  1341 => x"38bc9008",
  1342 => x"a007bc90",
  1343 => x"0c9d51a4",
  1344 => x"c02db5ac",
  1345 => x"08802e89",
  1346 => x"38bc9008",
  1347 => x"8107bc90",
  1348 => x"0c9b51a4",
  1349 => x"c02db5ac",
  1350 => x"08802e89",
  1351 => x"38bc9008",
  1352 => x"8207bc90",
  1353 => x"0c9c51a4",
  1354 => x"c02db5ac",
  1355 => x"08802e89",
  1356 => x"38bc9008",
  1357 => x"8407bc90",
  1358 => x"0ca351a4",
  1359 => x"c02db5ac",
  1360 => x"08802e89",
  1361 => x"38bc9008",
  1362 => x"8807bc90",
  1363 => x"0c81fd51",
  1364 => x"a4c02d81",
  1365 => x"fa51a4c0",
  1366 => x"2daf9704",
  1367 => x"81f551a4",
  1368 => x"c02db5ac",
  1369 => x"08812a70",
  1370 => x"81065152",
  1371 => x"71802eaf",
  1372 => x"38bc9c08",
  1373 => x"5271802e",
  1374 => x"8938ff12",
  1375 => x"bc9c0cab",
  1376 => x"9f04bc98",
  1377 => x"0810bc98",
  1378 => x"08057084",
  1379 => x"29165152",
  1380 => x"88120880",
  1381 => x"2e8938ff",
  1382 => x"51881208",
  1383 => x"52712d81",
  1384 => x"f251a4c0",
  1385 => x"2db5ac08",
  1386 => x"812a7081",
  1387 => x"06515271",
  1388 => x"802eb138",
  1389 => x"bc9808ff",
  1390 => x"11bc9c08",
  1391 => x"56535373",
  1392 => x"72258938",
  1393 => x"8114bc9c",
  1394 => x"0cabe404",
  1395 => x"72101370",
  1396 => x"84291651",
  1397 => x"52881208",
  1398 => x"802e8938",
  1399 => x"fe518812",
  1400 => x"0852712d",
  1401 => x"81fd51a4",
  1402 => x"c02db5ac",
  1403 => x"08812a70",
  1404 => x"81065152",
  1405 => x"71802e86",
  1406 => x"38800bbc",
  1407 => x"9c0c81fa",
  1408 => x"51a4c02d",
  1409 => x"b5ac0881",
  1410 => x"2a708106",
  1411 => x"51527180",
  1412 => x"2e8938bc",
  1413 => x"9808ff05",
  1414 => x"bc9c0cbc",
  1415 => x"9c087053",
  1416 => x"5473802e",
  1417 => x"8a388c15",
  1418 => x"ff155555",
  1419 => x"aca10482",
  1420 => x"0bb5c00c",
  1421 => x"718f06b5",
  1422 => x"bc0c81eb",
  1423 => x"51a4c02d",
  1424 => x"b5ac0881",
  1425 => x"2a708106",
  1426 => x"51527180",
  1427 => x"2ead3874",
  1428 => x"08852e09",
  1429 => x"8106a438",
  1430 => x"881580f5",
  1431 => x"2dff0552",
  1432 => x"71881681",
  1433 => x"b72d7198",
  1434 => x"2b527180",
  1435 => x"25883880",
  1436 => x"0b881681",
  1437 => x"b72d7451",
  1438 => x"a5b62d81",
  1439 => x"f451a4c0",
  1440 => x"2db5ac08",
  1441 => x"812a7081",
  1442 => x"06515271",
  1443 => x"802eb338",
  1444 => x"7408852e",
  1445 => x"098106aa",
  1446 => x"38881580",
  1447 => x"f52d8105",
  1448 => x"52718816",
  1449 => x"81b72d71",
  1450 => x"81ff068b",
  1451 => x"1680f52d",
  1452 => x"54527272",
  1453 => x"27873872",
  1454 => x"881681b7",
  1455 => x"2d7451a5",
  1456 => x"b62d80da",
  1457 => x"51a4c02d",
  1458 => x"b5ac0881",
  1459 => x"2a708106",
  1460 => x"51527180",
  1461 => x"2e80ff38",
  1462 => x"bc9408bc",
  1463 => x"9c085553",
  1464 => x"73802e8a",
  1465 => x"388c13ff",
  1466 => x"155553ad",
  1467 => x"e0047208",
  1468 => x"5271822e",
  1469 => x"a6387182",
  1470 => x"26893871",
  1471 => x"812ea938",
  1472 => x"aed60471",
  1473 => x"832eb138",
  1474 => x"71842e09",
  1475 => x"810680c6",
  1476 => x"38881308",
  1477 => x"51a7812d",
  1478 => x"aed604bc",
  1479 => x"9c085188",
  1480 => x"13085271",
  1481 => x"2daed604",
  1482 => x"810b8814",
  1483 => x"082bbc88",
  1484 => x"0832bc88",
  1485 => x"0caed304",
  1486 => x"881380f5",
  1487 => x"2d81058b",
  1488 => x"1480f52d",
  1489 => x"53547174",
  1490 => x"24833880",
  1491 => x"54738814",
  1492 => x"81b72da5",
  1493 => x"e62d8054",
  1494 => x"800bb5c0",
  1495 => x"0c738f06",
  1496 => x"b5bc0ca0",
  1497 => x"5273bc9c",
  1498 => x"082e0981",
  1499 => x"069838bc",
  1500 => x"9808ff05",
  1501 => x"74327009",
  1502 => x"81057072",
  1503 => x"079f2a91",
  1504 => x"71315151",
  1505 => x"53537151",
  1506 => x"82ee2d81",
  1507 => x"14548e74",
  1508 => x"25c638b5",
  1509 => x"a8085271",
  1510 => x"b5ac0c02",
  1511 => x"94050d04",
  1512 => x"00ffffff",
  1513 => x"ff00ffff",
  1514 => x"ffff00ff",
  1515 => x"ffffff00",
  1516 => x"52657365",
  1517 => x"74000000",
  1518 => x"53617665",
  1519 => x"20736574",
  1520 => x"74696e67",
  1521 => x"73000000",
  1522 => x"5363616e",
  1523 => x"6c696e65",
  1524 => x"73000000",
  1525 => x"4c6f6164",
  1526 => x"20524f4d",
  1527 => x"20100000",
  1528 => x"45786974",
  1529 => x"00000000",
  1530 => x"50432045",
  1531 => x"6e67696e",
  1532 => x"65206d6f",
  1533 => x"64650000",
  1534 => x"54757262",
  1535 => x"6f677261",
  1536 => x"66782031",
  1537 => x"36206d6f",
  1538 => x"64650000",
  1539 => x"56474120",
  1540 => x"2d203331",
  1541 => x"4b487a2c",
  1542 => x"20363048",
  1543 => x"7a000000",
  1544 => x"5456202d",
  1545 => x"20343830",
  1546 => x"692c2036",
  1547 => x"30487a00",
  1548 => x"4261636b",
  1549 => x"00000000",
  1550 => x"46504741",
  1551 => x"50434520",
  1552 => x"43464700",
  1553 => x"52656164",
  1554 => x"20666169",
  1555 => x"6c65640a",
  1556 => x"00000000",
  1557 => x"4661696c",
  1558 => x"65640a00",
  1559 => x"4c6f6164",
  1560 => x"696e6720",
  1561 => x"00000000",
  1562 => x"496e6974",
  1563 => x"69616c69",
  1564 => x"7a696e67",
  1565 => x"20534420",
  1566 => x"63617264",
  1567 => x"0a000000",
  1568 => x"424f4f54",
  1569 => x"20202020",
  1570 => x"50434500",
  1571 => x"43617264",
  1572 => x"20696e69",
  1573 => x"74206661",
  1574 => x"696c6564",
  1575 => x"0a000000",
  1576 => x"4d425220",
  1577 => x"6661696c",
  1578 => x"0a000000",
  1579 => x"46415431",
  1580 => x"36202020",
  1581 => x"00000000",
  1582 => x"46415433",
  1583 => x"32202020",
  1584 => x"00000000",
  1585 => x"4e6f2070",
  1586 => x"61727469",
  1587 => x"74696f6e",
  1588 => x"20736967",
  1589 => x"0a000000",
  1590 => x"42616420",
  1591 => x"70617274",
  1592 => x"0a000000",
  1593 => x"53444843",
  1594 => x"20657272",
  1595 => x"6f72210a",
  1596 => x"00000000",
  1597 => x"53442069",
  1598 => x"6e69742e",
  1599 => x"2e2e0a00",
  1600 => x"53442063",
  1601 => x"61726420",
  1602 => x"72657365",
  1603 => x"74206661",
  1604 => x"696c6564",
  1605 => x"210a0000",
  1606 => x"57726974",
  1607 => x"65206661",
  1608 => x"696c6564",
  1609 => x"0a000000",
  1610 => x"16200000",
  1611 => x"14200000",
  1612 => x"15200000",
  1613 => x"00000002",
  1614 => x"00000002",
  1615 => x"000017b0",
  1616 => x"000004ce",
  1617 => x"00000002",
  1618 => x"000017b8",
  1619 => x"000003a2",
  1620 => x"00000003",
  1621 => x"000019a0",
  1622 => x"00000002",
  1623 => x"00000001",
  1624 => x"000017c8",
  1625 => x"00000001",
  1626 => x"00000003",
  1627 => x"00001998",
  1628 => x"00000002",
  1629 => x"00000002",
  1630 => x"000017d4",
  1631 => x"0000062e",
  1632 => x"00000002",
  1633 => x"000017e0",
  1634 => x"000012a3",
  1635 => x"00000000",
  1636 => x"00000000",
  1637 => x"00000000",
  1638 => x"000017e8",
  1639 => x"000017f8",
  1640 => x"0000180c",
  1641 => x"00001820",
  1642 => x"00000002",
  1643 => x"00001ad8",
  1644 => x"000004e3",
  1645 => x"00000002",
  1646 => x"00001ae8",
  1647 => x"000004e3",
  1648 => x"00000002",
  1649 => x"00001af8",
  1650 => x"000004e3",
  1651 => x"00000002",
  1652 => x"00001b08",
  1653 => x"000004e3",
  1654 => x"00000002",
  1655 => x"00001b18",
  1656 => x"000004e3",
  1657 => x"00000002",
  1658 => x"00001b28",
  1659 => x"000004e3",
  1660 => x"00000002",
  1661 => x"00001b38",
  1662 => x"000004e3",
  1663 => x"00000002",
  1664 => x"00001b48",
  1665 => x"000004e3",
  1666 => x"00000002",
  1667 => x"00001b58",
  1668 => x"000004e3",
  1669 => x"00000002",
  1670 => x"00001b68",
  1671 => x"000004e3",
  1672 => x"00000002",
  1673 => x"00001b78",
  1674 => x"000004e3",
  1675 => x"00000002",
  1676 => x"00001b88",
  1677 => x"000004e3",
  1678 => x"00000002",
  1679 => x"00001b98",
  1680 => x"000004e3",
  1681 => x"00000004",
  1682 => x"00001830",
  1683 => x"00001938",
  1684 => x"00000000",
  1685 => x"00000000",
  1686 => x"000005c2",
  1687 => x"00000000",
  1688 => x"00000000",
  1689 => x"00000000",
  1690 => x"00000000",
  1691 => x"00000000",
  1692 => x"00000000",
  1693 => x"00000000",
  1694 => x"00000000",
  1695 => x"00000000",
  1696 => x"00000000",
  1697 => x"00000000",
  1698 => x"00000000",
  1699 => x"00000000",
  1700 => x"00000000",
  1701 => x"00000000",
  1702 => x"00000000",
  1703 => x"00000000",
  1704 => x"00000000",
  1705 => x"00000000",
  1706 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

