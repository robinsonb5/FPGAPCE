-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb0",
     9 => x"d0080b0b",
    10 => x"0bb0d408",
    11 => x"0b0b0bb0",
    12 => x"d8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b0d80c0b",
    16 => x"0b0bb0d4",
    17 => x"0c0b0b0b",
    18 => x"b0d00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0baa98",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b0d070b7",
    57 => x"bc278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8b970402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b0e00c9f",
    65 => x"0bb0e40c",
    66 => x"a0717081",
    67 => x"055334b0",
    68 => x"e408ff05",
    69 => x"b0e40cb0",
    70 => x"e4088025",
    71 => x"eb38b0e0",
    72 => x"08ff05b0",
    73 => x"e00cb0e0",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb0e0",
    94 => x"08258f38",
    95 => x"82b22db0",
    96 => x"e008ff05",
    97 => x"b0e00c82",
    98 => x"f404b0e0",
    99 => x"08b0e408",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b0e008",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b0",
   108 => x"e4088105",
   109 => x"b0e40cb0",
   110 => x"e408519f",
   111 => x"7125e238",
   112 => x"800bb0e4",
   113 => x"0cb0e008",
   114 => x"8105b0e0",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b0e40881",
   120 => x"05b0e40c",
   121 => x"b0e408a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b0e40cb0",
   125 => x"e0088105",
   126 => x"b0e00c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb0",
   155 => x"e80cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb0e8",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b0e80884",
   167 => x"07b0e80c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0bad",
   172 => x"dc0c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cb0e808",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f4050d",
   198 => x"74708206",
   199 => x"b7ac0cad",
   200 => x"f8718106",
   201 => x"54545171",
   202 => x"881481b7",
   203 => x"2d70822a",
   204 => x"70810651",
   205 => x"51709414",
   206 => x"81b72d70",
   207 => x"b0d00c02",
   208 => x"8c050d04",
   209 => x"02f4050d",
   210 => x"abb052b0",
   211 => x"f05194a2",
   212 => x"2db0d008",
   213 => x"802e9538",
   214 => x"b2cc52b0",
   215 => x"f05196d8",
   216 => x"2db2cc08",
   217 => x"70fec00c",
   218 => x"5186942d",
   219 => x"028c050d",
   220 => x"0402f805",
   221 => x"0db7ac08",
   222 => x"8206ae80",
   223 => x"0b80f52d",
   224 => x"52527080",
   225 => x"2e853871",
   226 => x"810752ae",
   227 => x"8c0b80f5",
   228 => x"2d517080",
   229 => x"2e853871",
   230 => x"84075271",
   231 => x"b0d00c02",
   232 => x"88050d04",
   233 => x"02f0050d",
   234 => x"86f12db0",
   235 => x"d008abb0",
   236 => x"53b0f052",
   237 => x"5394a22d",
   238 => x"b0d00880",
   239 => x"2ea33872",
   240 => x"b2cc0cb2",
   241 => x"d05480fd",
   242 => x"53807470",
   243 => x"8405560c",
   244 => x"ff135372",
   245 => x"8025f238",
   246 => x"b2cc52b0",
   247 => x"f05196fe",
   248 => x"2d029005",
   249 => x"0d0402d8",
   250 => x"050d810b",
   251 => x"fec40c84",
   252 => x"0bfec40c",
   253 => x"7b52b0f0",
   254 => x"5194a22d",
   255 => x"b0d00853",
   256 => x"b0d00880",
   257 => x"2e81c038",
   258 => x"abbc5185",
   259 => x"f32db0f4",
   260 => x"0856800b",
   261 => x"ff175859",
   262 => x"76792e8b",
   263 => x"38811977",
   264 => x"812a5859",
   265 => x"76f738f7",
   266 => x"19769fff",
   267 => x"06545972",
   268 => x"802e8b38",
   269 => x"fc8016b0",
   270 => x"f0525696",
   271 => x"ab2d8076",
   272 => x"2580fd38",
   273 => x"78527651",
   274 => x"84802db2",
   275 => x"cc52b0f0",
   276 => x"5196d82d",
   277 => x"b0d00853",
   278 => x"b0d00880",
   279 => x"2e80c838",
   280 => x"b2cc5a80",
   281 => x"58899404",
   282 => x"79708405",
   283 => x"5b087083",
   284 => x"fe800671",
   285 => x"882b83fe",
   286 => x"80067188",
   287 => x"2a077288",
   288 => x"2a83fe80",
   289 => x"0673982a",
   290 => x"07fec80c",
   291 => x"fec80c56",
   292 => x"84195953",
   293 => x"75538480",
   294 => x"76258438",
   295 => x"84805372",
   296 => x"7824c538",
   297 => x"89b004ab",
   298 => x"cc5185f3",
   299 => x"2d89c704",
   300 => x"b0f05196",
   301 => x"ab2dfc80",
   302 => x"16811858",
   303 => x"5688be04",
   304 => x"820bfec4",
   305 => x"0c815372",
   306 => x"b0d00c02",
   307 => x"a8050d04",
   308 => x"a3d42d04",
   309 => x"02ec050d",
   310 => x"81175480",
   311 => x"5573752e",
   312 => x"a3387451",
   313 => x"93cd2db0",
   314 => x"d008b0d0",
   315 => x"08098105",
   316 => x"70b0d008",
   317 => x"079f2a76",
   318 => x"71318119",
   319 => x"59575153",
   320 => x"5373df38",
   321 => x"72802e98",
   322 => x"38800b8b",
   323 => x"1481b72d",
   324 => x"abdc5185",
   325 => x"f32d7251",
   326 => x"85f32d72",
   327 => x"5187e62d",
   328 => x"ade051a5",
   329 => x"b22da3d4",
   330 => x"2d805184",
   331 => x"e52d0294",
   332 => x"050d0402",
   333 => x"e8050d80",
   334 => x"705755b6",
   335 => x"d808752e",
   336 => x"80ca3874",
   337 => x"5193cd2d",
   338 => x"b0d00880",
   339 => x"2eae3875",
   340 => x"9029b0fc",
   341 => x"058117b0",
   342 => x"d0085657",
   343 => x"528a5373",
   344 => x"70810555",
   345 => x"80f52d72",
   346 => x"70810554",
   347 => x"81b72dff",
   348 => x"13537280",
   349 => x"25e93880",
   350 => x"7281b72d",
   351 => x"81155575",
   352 => x"8b248938",
   353 => x"b6d80875",
   354 => x"26ffb838",
   355 => x"aed051a5",
   356 => x"b22d0298",
   357 => x"050d0402",
   358 => x"f4050d80",
   359 => x"5186942d",
   360 => x"810bfec4",
   361 => x"0c800bfe",
   362 => x"c00c840b",
   363 => x"fec40c83",
   364 => x"0bfecc0c",
   365 => x"a1b52da3",
   366 => x"c82da19a",
   367 => x"2da19a2d",
   368 => x"81f72d81",
   369 => x"5184e52d",
   370 => x"a19a2da1",
   371 => x"9a2d8151",
   372 => x"84e52dab",
   373 => x"e85185f3",
   374 => x"2d9bb12d",
   375 => x"b0d00880",
   376 => x"2e818938",
   377 => x"8dbb2db0",
   378 => x"d00852b0",
   379 => x"d0088a38",
   380 => x"ac805185",
   381 => x"f32d8cf4",
   382 => x"0486c42d",
   383 => x"ac945187",
   384 => x"e62db0d0",
   385 => x"08802e89",
   386 => x"38805184",
   387 => x"e52d8c97",
   388 => x"04aca051",
   389 => x"85f32dad",
   390 => x"e051a5b2",
   391 => x"2da1cd2d",
   392 => x"a5c22db0",
   393 => x"d0085386",
   394 => x"f12db0d0",
   395 => x"08fec00c",
   396 => x"86f12db0",
   397 => x"d008b0ec",
   398 => x"082e9c38",
   399 => x"b0d008b0",
   400 => x"ec0c8452",
   401 => x"725184e5",
   402 => x"2da19a2d",
   403 => x"a19a2dff",
   404 => x"12527180",
   405 => x"25ee3872",
   406 => x"802e8938",
   407 => x"8a0bfec4",
   408 => x"0c8c9d04",
   409 => x"820bfec4",
   410 => x"0c8c9d04",
   411 => x"acb45185",
   412 => x"f32d8052",
   413 => x"71b0d00c",
   414 => x"028c050d",
   415 => x"0402e805",
   416 => x"0d77797b",
   417 => x"58555580",
   418 => x"53727625",
   419 => x"a3387470",
   420 => x"81055680",
   421 => x"f52d7470",
   422 => x"81055680",
   423 => x"f52d5252",
   424 => x"71712e86",
   425 => x"3881518d",
   426 => x"b2048113",
   427 => x"538d8904",
   428 => x"805170b0",
   429 => x"d00c0298",
   430 => x"050d0402",
   431 => x"d8050d80",
   432 => x"0bb6d40c",
   433 => x"b2cc5280",
   434 => x"519e992d",
   435 => x"b0d00854",
   436 => x"b0d0088c",
   437 => x"38acc851",
   438 => x"85f32d73",
   439 => x"5592d604",
   440 => x"8056810b",
   441 => x"b6f80c88",
   442 => x"53acd452",
   443 => x"b382518c",
   444 => x"fd2db0d0",
   445 => x"08762e09",
   446 => x"81068738",
   447 => x"b0d008b6",
   448 => x"f80c8853",
   449 => x"ace052b3",
   450 => x"9e518cfd",
   451 => x"2db0d008",
   452 => x"8738b0d0",
   453 => x"08b6f80c",
   454 => x"b6f80880",
   455 => x"2e80f638",
   456 => x"b6920b80",
   457 => x"f52db693",
   458 => x"0b80f52d",
   459 => x"71982b71",
   460 => x"902b07b6",
   461 => x"940b80f5",
   462 => x"2d70882b",
   463 => x"7207b695",
   464 => x"0b80f52d",
   465 => x"7107b6ca",
   466 => x"0b80f52d",
   467 => x"b6cb0b80",
   468 => x"f52d7188",
   469 => x"2b07535f",
   470 => x"54525a56",
   471 => x"57557381",
   472 => x"abaa2e09",
   473 => x"81068d38",
   474 => x"75519fb4",
   475 => x"2db0d008",
   476 => x"568f8104",
   477 => x"7382d4d5",
   478 => x"2e8738ac",
   479 => x"ec518fc2",
   480 => x"04b2cc52",
   481 => x"75519e99",
   482 => x"2db0d008",
   483 => x"55b0d008",
   484 => x"802e83c2",
   485 => x"388853ac",
   486 => x"e052b39e",
   487 => x"518cfd2d",
   488 => x"b0d00889",
   489 => x"38810bb6",
   490 => x"d40c8fc8",
   491 => x"048853ac",
   492 => x"d452b382",
   493 => x"518cfd2d",
   494 => x"b0d00880",
   495 => x"2e8a38ad",
   496 => x"805185f3",
   497 => x"2d90a204",
   498 => x"b6ca0b80",
   499 => x"f52d5473",
   500 => x"80d52e09",
   501 => x"810680ca",
   502 => x"38b6cb0b",
   503 => x"80f52d54",
   504 => x"7381aa2e",
   505 => x"098106ba",
   506 => x"38800bb2",
   507 => x"cc0b80f5",
   508 => x"2d565474",
   509 => x"81e92e83",
   510 => x"38815474",
   511 => x"81eb2e8c",
   512 => x"38805573",
   513 => x"752e0981",
   514 => x"0682cb38",
   515 => x"b2d70b80",
   516 => x"f52d5574",
   517 => x"8d38b2d8",
   518 => x"0b80f52d",
   519 => x"5473822e",
   520 => x"86388055",
   521 => x"92d604b2",
   522 => x"d90b80f5",
   523 => x"2d70b6cc",
   524 => x"0cff05b6",
   525 => x"d00cb2da",
   526 => x"0b80f52d",
   527 => x"b2db0b80",
   528 => x"f52d5876",
   529 => x"05778280",
   530 => x"290570b6",
   531 => x"dc0cb2dc",
   532 => x"0b80f52d",
   533 => x"70b6f00c",
   534 => x"b6d40859",
   535 => x"57587680",
   536 => x"2e81a338",
   537 => x"8853ace0",
   538 => x"52b39e51",
   539 => x"8cfd2db0",
   540 => x"d00881e2",
   541 => x"38b6cc08",
   542 => x"70842bb6",
   543 => x"d80c70b6",
   544 => x"ec0cb2f1",
   545 => x"0b80f52d",
   546 => x"b2f00b80",
   547 => x"f52d7182",
   548 => x"802905b2",
   549 => x"f20b80f5",
   550 => x"2d708480",
   551 => x"802912b2",
   552 => x"f30b80f5",
   553 => x"2d708180",
   554 => x"0a291270",
   555 => x"b6f40cb6",
   556 => x"f0087129",
   557 => x"b6dc0805",
   558 => x"70b6e00c",
   559 => x"b2f90b80",
   560 => x"f52db2f8",
   561 => x"0b80f52d",
   562 => x"71828029",
   563 => x"05b2fa0b",
   564 => x"80f52d70",
   565 => x"84808029",
   566 => x"12b2fb0b",
   567 => x"80f52d70",
   568 => x"982b81f0",
   569 => x"0a067205",
   570 => x"70b6e40c",
   571 => x"fe117e29",
   572 => x"7705b6e8",
   573 => x"0c525952",
   574 => x"43545e51",
   575 => x"5259525d",
   576 => x"57595792",
   577 => x"d404b2de",
   578 => x"0b80f52d",
   579 => x"b2dd0b80",
   580 => x"f52d7182",
   581 => x"80290570",
   582 => x"b6d80c70",
   583 => x"a02983ff",
   584 => x"0570892a",
   585 => x"70b6ec0c",
   586 => x"b2e30b80",
   587 => x"f52db2e2",
   588 => x"0b80f52d",
   589 => x"71828029",
   590 => x"0570b6f4",
   591 => x"0c7b7129",
   592 => x"1e70b6e8",
   593 => x"0c7db6e4",
   594 => x"0c7305b6",
   595 => x"e00c555e",
   596 => x"51515555",
   597 => x"815574b0",
   598 => x"d00c02a8",
   599 => x"050d0402",
   600 => x"ec050d76",
   601 => x"70872c71",
   602 => x"80ff0655",
   603 => x"5654b6d4",
   604 => x"088a3873",
   605 => x"882c7481",
   606 => x"ff065455",
   607 => x"b2cc52b6",
   608 => x"dc081551",
   609 => x"9e992db0",
   610 => x"d00854b0",
   611 => x"d008802e",
   612 => x"b338b6d4",
   613 => x"08802e98",
   614 => x"38728429",
   615 => x"b2cc0570",
   616 => x"0852539f",
   617 => x"b42db0d0",
   618 => x"08f00a06",
   619 => x"5393c204",
   620 => x"7210b2cc",
   621 => x"057080e0",
   622 => x"2d52539f",
   623 => x"e42db0d0",
   624 => x"08537254",
   625 => x"73b0d00c",
   626 => x"0294050d",
   627 => x"0402ec05",
   628 => x"0d767084",
   629 => x"2cb6e808",
   630 => x"05718f06",
   631 => x"52555372",
   632 => x"8938b2cc",
   633 => x"5273519e",
   634 => x"992d72a0",
   635 => x"29b2cc05",
   636 => x"54807480",
   637 => x"f52d5455",
   638 => x"72752e83",
   639 => x"38815572",
   640 => x"81e52e93",
   641 => x"3874802e",
   642 => x"8e388b14",
   643 => x"80f52d98",
   644 => x"06537280",
   645 => x"2e833880",
   646 => x"5473b0d0",
   647 => x"0c029405",
   648 => x"0d0402cc",
   649 => x"050d7e60",
   650 => x"5e5a800b",
   651 => x"b6e408b6",
   652 => x"e808595c",
   653 => x"568058b6",
   654 => x"d808782e",
   655 => x"81ae3877",
   656 => x"8f06a017",
   657 => x"5754738f",
   658 => x"38b2cc52",
   659 => x"76518117",
   660 => x"579e992d",
   661 => x"b2cc5680",
   662 => x"7680f52d",
   663 => x"56547474",
   664 => x"2e833881",
   665 => x"547481e5",
   666 => x"2e80f638",
   667 => x"81707506",
   668 => x"555c7380",
   669 => x"2e80ea38",
   670 => x"8b1680f5",
   671 => x"2d980659",
   672 => x"7880de38",
   673 => x"8b537c52",
   674 => x"75518cfd",
   675 => x"2db0d008",
   676 => x"80cf389c",
   677 => x"1608519f",
   678 => x"b42db0d0",
   679 => x"08841b0c",
   680 => x"9a1680e0",
   681 => x"2d519fe4",
   682 => x"2db0d008",
   683 => x"b0d00888",
   684 => x"1c0cb0d0",
   685 => x"085555b6",
   686 => x"d408802e",
   687 => x"98389416",
   688 => x"80e02d51",
   689 => x"9fe42db0",
   690 => x"d008902b",
   691 => x"83fff00a",
   692 => x"06701651",
   693 => x"5473881b",
   694 => x"0c787a0c",
   695 => x"7b5496a2",
   696 => x"04811858",
   697 => x"b6d80878",
   698 => x"26fed438",
   699 => x"b6d40880",
   700 => x"2eae387a",
   701 => x"5192df2d",
   702 => x"b0d008b0",
   703 => x"d00880ff",
   704 => x"fffff806",
   705 => x"555b7380",
   706 => x"fffffff8",
   707 => x"2e9238b0",
   708 => x"d008fe05",
   709 => x"b6cc0829",
   710 => x"b6e00805",
   711 => x"5794b504",
   712 => x"805473b0",
   713 => x"d00c02b4",
   714 => x"050d0402",
   715 => x"f4050d74",
   716 => x"70088105",
   717 => x"710c7008",
   718 => x"b6d00806",
   719 => x"5353718e",
   720 => x"38881308",
   721 => x"5192df2d",
   722 => x"b0d00888",
   723 => x"140c810b",
   724 => x"b0d00c02",
   725 => x"8c050d04",
   726 => x"02f0050d",
   727 => x"75881108",
   728 => x"fe05b6cc",
   729 => x"0829b6e0",
   730 => x"08117208",
   731 => x"b6d00806",
   732 => x"05795553",
   733 => x"54549e99",
   734 => x"2d029005",
   735 => x"0d0402f0",
   736 => x"050d7588",
   737 => x"1108fe05",
   738 => x"b6cc0829",
   739 => x"b6e00811",
   740 => x"7208b6d0",
   741 => x"08060579",
   742 => x"55535454",
   743 => x"9cd92d02",
   744 => x"90050d04",
   745 => x"02f4050d",
   746 => x"d45281ff",
   747 => x"720c7108",
   748 => x"5381ff72",
   749 => x"0c72882b",
   750 => x"83fe8006",
   751 => x"72087081",
   752 => x"ff065152",
   753 => x"5381ff72",
   754 => x"0c727107",
   755 => x"882b7208",
   756 => x"7081ff06",
   757 => x"51525381",
   758 => x"ff720c72",
   759 => x"7107882b",
   760 => x"72087081",
   761 => x"ff067207",
   762 => x"b0d00c52",
   763 => x"53028c05",
   764 => x"0d0402f4",
   765 => x"050d7476",
   766 => x"7181ff06",
   767 => x"d40c5353",
   768 => x"b6fc0885",
   769 => x"3871892b",
   770 => x"5271982a",
   771 => x"d40c7190",
   772 => x"2a7081ff",
   773 => x"06d40c51",
   774 => x"71882a70",
   775 => x"81ff06d4",
   776 => x"0c517181",
   777 => x"ff06d40c",
   778 => x"72902a70",
   779 => x"81ff06d4",
   780 => x"0c51d408",
   781 => x"7081ff06",
   782 => x"515182b8",
   783 => x"bf527081",
   784 => x"ff2e0981",
   785 => x"06943881",
   786 => x"ff0bd40c",
   787 => x"d4087081",
   788 => x"ff06ff14",
   789 => x"54515171",
   790 => x"e53870b0",
   791 => x"d00c028c",
   792 => x"050d0402",
   793 => x"fc050d81",
   794 => x"c75181ff",
   795 => x"0bd40cff",
   796 => x"11517080",
   797 => x"25f43802",
   798 => x"84050d04",
   799 => x"02f0050d",
   800 => x"98e32d8f",
   801 => x"cf538052",
   802 => x"87fc80f7",
   803 => x"5197f22d",
   804 => x"b0d00854",
   805 => x"b0d00881",
   806 => x"2e098106",
   807 => x"a33881ff",
   808 => x"0bd40c82",
   809 => x"0a52849c",
   810 => x"80e95197",
   811 => x"f22db0d0",
   812 => x"088b3881",
   813 => x"ff0bd40c",
   814 => x"735399c6",
   815 => x"0498e32d",
   816 => x"ff135372",
   817 => x"c13872b0",
   818 => x"d00c0290",
   819 => x"050d0402",
   820 => x"f4050d81",
   821 => x"ff0bd40c",
   822 => x"93538052",
   823 => x"87fc80c1",
   824 => x"5197f22d",
   825 => x"b0d0088b",
   826 => x"3881ff0b",
   827 => x"d40c8153",
   828 => x"99fc0498",
   829 => x"e32dff13",
   830 => x"5372df38",
   831 => x"72b0d00c",
   832 => x"028c050d",
   833 => x"0402f005",
   834 => x"0d98e32d",
   835 => x"83aa5284",
   836 => x"9c80c851",
   837 => x"97f22db0",
   838 => x"d008812e",
   839 => x"09810692",
   840 => x"3897a42d",
   841 => x"b0d00883",
   842 => x"ffff0653",
   843 => x"7283aa2e",
   844 => x"973899cf",
   845 => x"2d9ac304",
   846 => x"81549ba8",
   847 => x"04ad8c51",
   848 => x"85f32d80",
   849 => x"549ba804",
   850 => x"81ff0bd4",
   851 => x"0cb15398",
   852 => x"fc2db0d0",
   853 => x"08802e80",
   854 => x"c0388052",
   855 => x"87fc80fa",
   856 => x"5197f22d",
   857 => x"b0d008b1",
   858 => x"3881ff0b",
   859 => x"d40cd408",
   860 => x"5381ff0b",
   861 => x"d40c81ff",
   862 => x"0bd40c81",
   863 => x"ff0bd40c",
   864 => x"81ff0bd4",
   865 => x"0c72862a",
   866 => x"708106b0",
   867 => x"d0085651",
   868 => x"5372802e",
   869 => x"93389ab8",
   870 => x"0472822e",
   871 => x"ff9f38ff",
   872 => x"135372ff",
   873 => x"aa387254",
   874 => x"73b0d00c",
   875 => x"0290050d",
   876 => x"0402f005",
   877 => x"0d810bb6",
   878 => x"fc0c8454",
   879 => x"d008708f",
   880 => x"2a708106",
   881 => x"51515372",
   882 => x"f33872d0",
   883 => x"0c98e32d",
   884 => x"ad9c5185",
   885 => x"f32dd008",
   886 => x"708f2a70",
   887 => x"81065151",
   888 => x"5372f338",
   889 => x"810bd00c",
   890 => x"b1538052",
   891 => x"84d480c0",
   892 => x"5197f22d",
   893 => x"b0d00881",
   894 => x"2ea13872",
   895 => x"822e0981",
   896 => x"068c38ad",
   897 => x"a85185f3",
   898 => x"2d80539c",
   899 => x"d004ff13",
   900 => x"5372d738",
   901 => x"ff145473",
   902 => x"ffa2389a",
   903 => x"852db0d0",
   904 => x"08b6fc0c",
   905 => x"b0d0088b",
   906 => x"38815287",
   907 => x"fc80d051",
   908 => x"97f22d81",
   909 => x"ff0bd40c",
   910 => x"d008708f",
   911 => x"2a708106",
   912 => x"51515372",
   913 => x"f33872d0",
   914 => x"0c81ff0b",
   915 => x"d40c8153",
   916 => x"72b0d00c",
   917 => x"0290050d",
   918 => x"0402e805",
   919 => x"0d785681",
   920 => x"ff0bd40c",
   921 => x"d008708f",
   922 => x"2a708106",
   923 => x"51515372",
   924 => x"f3388281",
   925 => x"0bd00c81",
   926 => x"ff0bd40c",
   927 => x"775287fc",
   928 => x"80d85197",
   929 => x"f22db0d0",
   930 => x"08802e8c",
   931 => x"38adc051",
   932 => x"85f32d81",
   933 => x"539e9004",
   934 => x"81ff0bd4",
   935 => x"0c81fe0b",
   936 => x"d40c80ff",
   937 => x"55757084",
   938 => x"05570870",
   939 => x"982ad40c",
   940 => x"70902c70",
   941 => x"81ff06d4",
   942 => x"0c547088",
   943 => x"2c7081ff",
   944 => x"06d40c54",
   945 => x"7081ff06",
   946 => x"d40c54ff",
   947 => x"15557480",
   948 => x"25d33881",
   949 => x"ff0bd40c",
   950 => x"81ff0bd4",
   951 => x"0c81ff0b",
   952 => x"d40c868d",
   953 => x"a05481ff",
   954 => x"0bd40cd4",
   955 => x"0881ff06",
   956 => x"55748738",
   957 => x"ff145473",
   958 => x"ed3881ff",
   959 => x"0bd40cd0",
   960 => x"08708f2a",
   961 => x"70810651",
   962 => x"515372f3",
   963 => x"3872d00c",
   964 => x"72b0d00c",
   965 => x"0298050d",
   966 => x"0402e805",
   967 => x"0d785580",
   968 => x"5681ff0b",
   969 => x"d40cd008",
   970 => x"708f2a70",
   971 => x"81065151",
   972 => x"5372f338",
   973 => x"82810bd0",
   974 => x"0c81ff0b",
   975 => x"d40c7752",
   976 => x"87fc80d1",
   977 => x"5197f22d",
   978 => x"80dbc6df",
   979 => x"54b0d008",
   980 => x"802e8a38",
   981 => x"abcc5185",
   982 => x"f32d9fab",
   983 => x"0481ff0b",
   984 => x"d40cd408",
   985 => x"7081ff06",
   986 => x"51537281",
   987 => x"fe2e0981",
   988 => x"069d3880",
   989 => x"ff5397a4",
   990 => x"2db0d008",
   991 => x"75708405",
   992 => x"570cff13",
   993 => x"53728025",
   994 => x"ed388156",
   995 => x"9f9504ff",
   996 => x"145473c9",
   997 => x"3881ff0b",
   998 => x"d40cd008",
   999 => x"708f2a70",
  1000 => x"81065151",
  1001 => x"5372f338",
  1002 => x"72d00c75",
  1003 => x"b0d00c02",
  1004 => x"98050d04",
  1005 => x"02f4050d",
  1006 => x"7470882a",
  1007 => x"83fe8006",
  1008 => x"7072982a",
  1009 => x"0772882b",
  1010 => x"87fc8080",
  1011 => x"0673982b",
  1012 => x"81f00a06",
  1013 => x"71730707",
  1014 => x"b0d00c56",
  1015 => x"51535102",
  1016 => x"8c050d04",
  1017 => x"02f8050d",
  1018 => x"028e0580",
  1019 => x"f52d7488",
  1020 => x"2b077083",
  1021 => x"ffff06b0",
  1022 => x"d00c5102",
  1023 => x"88050d04",
  1024 => x"02fc050d",
  1025 => x"72518071",
  1026 => x"0c800b84",
  1027 => x"120c0284",
  1028 => x"050d0402",
  1029 => x"f0050d75",
  1030 => x"70088412",
  1031 => x"08535353",
  1032 => x"ff547171",
  1033 => x"2ea838a3",
  1034 => x"ce2d8413",
  1035 => x"08708429",
  1036 => x"14881170",
  1037 => x"087081ff",
  1038 => x"06841808",
  1039 => x"81118706",
  1040 => x"841a0c53",
  1041 => x"51555151",
  1042 => x"51a3c82d",
  1043 => x"715473b0",
  1044 => x"d00c0290",
  1045 => x"050d0402",
  1046 => x"f8050da3",
  1047 => x"ce2de008",
  1048 => x"708b2a70",
  1049 => x"81065152",
  1050 => x"5270802e",
  1051 => x"9d38b780",
  1052 => x"08708429",
  1053 => x"b7880573",
  1054 => x"81ff0671",
  1055 => x"0c5151b7",
  1056 => x"80088111",
  1057 => x"8706b780",
  1058 => x"0c51800b",
  1059 => x"b7a80ca3",
  1060 => x"c12da3c8",
  1061 => x"2d028805",
  1062 => x"0d0402fc",
  1063 => x"050da3ce",
  1064 => x"2d810bb7",
  1065 => x"a80ca3c8",
  1066 => x"2db7a808",
  1067 => x"5170fa38",
  1068 => x"0284050d",
  1069 => x"0402fc05",
  1070 => x"0db78051",
  1071 => x"a0802da0",
  1072 => x"d751a3bd",
  1073 => x"2da2e72d",
  1074 => x"0284050d",
  1075 => x"0402f405",
  1076 => x"0da2cf04",
  1077 => x"b0d00881",
  1078 => x"f02e0981",
  1079 => x"06893881",
  1080 => x"0bb0c40c",
  1081 => x"a2cf04b0",
  1082 => x"d00881e0",
  1083 => x"2e098106",
  1084 => x"8938810b",
  1085 => x"b0c80ca2",
  1086 => x"cf04b0d0",
  1087 => x"0852b0c8",
  1088 => x"08802e88",
  1089 => x"38b0d008",
  1090 => x"81800552",
  1091 => x"71842c72",
  1092 => x"8f065353",
  1093 => x"b0c40880",
  1094 => x"2e993872",
  1095 => x"8429b084",
  1096 => x"05721381",
  1097 => x"712b7009",
  1098 => x"73080673",
  1099 => x"0c515353",
  1100 => x"a2c50472",
  1101 => x"8429b084",
  1102 => x"05721383",
  1103 => x"712b7208",
  1104 => x"07720c53",
  1105 => x"53800bb0",
  1106 => x"c80c800b",
  1107 => x"b0c40cb7",
  1108 => x"8051a093",
  1109 => x"2db0d008",
  1110 => x"ff24fef8",
  1111 => x"38800bb0",
  1112 => x"d00c028c",
  1113 => x"050d0402",
  1114 => x"f8050db0",
  1115 => x"84528f51",
  1116 => x"80727084",
  1117 => x"05540cff",
  1118 => x"11517080",
  1119 => x"25f23802",
  1120 => x"88050d04",
  1121 => x"02f0050d",
  1122 => x"7551a3ce",
  1123 => x"2d70822c",
  1124 => x"fc06b084",
  1125 => x"1172109e",
  1126 => x"06710870",
  1127 => x"722a7083",
  1128 => x"0682742b",
  1129 => x"70097406",
  1130 => x"760c5451",
  1131 => x"56575351",
  1132 => x"53a3c82d",
  1133 => x"71b0d00c",
  1134 => x"0290050d",
  1135 => x"0471980c",
  1136 => x"04ffb008",
  1137 => x"b0d00c04",
  1138 => x"810bffb0",
  1139 => x"0c04800b",
  1140 => x"ffb00c04",
  1141 => x"02fc050d",
  1142 => x"800bb0cc",
  1143 => x"0c805184",
  1144 => x"e52d0284",
  1145 => x"050d0402",
  1146 => x"ec050d76",
  1147 => x"54805287",
  1148 => x"0b881580",
  1149 => x"f52d5653",
  1150 => x"74722483",
  1151 => x"38a05372",
  1152 => x"5182ee2d",
  1153 => x"81128b15",
  1154 => x"80f52d54",
  1155 => x"52727225",
  1156 => x"de380294",
  1157 => x"050d0402",
  1158 => x"f0050db7",
  1159 => x"b0085481",
  1160 => x"f72d800b",
  1161 => x"b7b40c73",
  1162 => x"08802e81",
  1163 => x"8038820b",
  1164 => x"b0e40cb7",
  1165 => x"b4088f06",
  1166 => x"b0e00c73",
  1167 => x"08527183",
  1168 => x"2e963871",
  1169 => x"83268938",
  1170 => x"71812eaf",
  1171 => x"38a59804",
  1172 => x"71852e9f",
  1173 => x"38a59804",
  1174 => x"881480f5",
  1175 => x"2d841508",
  1176 => x"add05354",
  1177 => x"5285f32d",
  1178 => x"71842913",
  1179 => x"70085252",
  1180 => x"a59c0473",
  1181 => x"51a3e72d",
  1182 => x"a59804b7",
  1183 => x"ac088815",
  1184 => x"082c7081",
  1185 => x"06515271",
  1186 => x"802e8738",
  1187 => x"add451a5",
  1188 => x"9504add8",
  1189 => x"5185f32d",
  1190 => x"84140851",
  1191 => x"85f32db7",
  1192 => x"b4088105",
  1193 => x"b7b40c8c",
  1194 => x"1454a4a7",
  1195 => x"04029005",
  1196 => x"0d0471b7",
  1197 => x"b00ca497",
  1198 => x"2db7b408",
  1199 => x"ff05b7b8",
  1200 => x"0c0402ec",
  1201 => x"050db7b0",
  1202 => x"085580f8",
  1203 => x"51a3842d",
  1204 => x"b0d00881",
  1205 => x"2a708106",
  1206 => x"5152719b",
  1207 => x"388751a3",
  1208 => x"842db0d0",
  1209 => x"08812a70",
  1210 => x"81065152",
  1211 => x"71802eb1",
  1212 => x"38a5f704",
  1213 => x"a1cd2d87",
  1214 => x"51a3842d",
  1215 => x"b0d008f4",
  1216 => x"38a68704",
  1217 => x"a1cd2d80",
  1218 => x"f851a384",
  1219 => x"2db0d008",
  1220 => x"f338b0cc",
  1221 => x"08813270",
  1222 => x"b0cc0c70",
  1223 => x"525284e5",
  1224 => x"2db0cc08",
  1225 => x"a23880da",
  1226 => x"51a3842d",
  1227 => x"81f551a3",
  1228 => x"842d81f2",
  1229 => x"51a3842d",
  1230 => x"81eb51a3",
  1231 => x"842d81f4",
  1232 => x"51a3842d",
  1233 => x"aa8f0481",
  1234 => x"f551a384",
  1235 => x"2db0d008",
  1236 => x"812a7081",
  1237 => x"06515271",
  1238 => x"802e8f38",
  1239 => x"b7b80852",
  1240 => x"71802e86",
  1241 => x"38ff12b7",
  1242 => x"b80c81f2",
  1243 => x"51a3842d",
  1244 => x"b0d00881",
  1245 => x"2a708106",
  1246 => x"51527180",
  1247 => x"2e9538b7",
  1248 => x"b408ff05",
  1249 => x"b7b80854",
  1250 => x"52727225",
  1251 => x"86388113",
  1252 => x"b7b80cb7",
  1253 => x"b8087053",
  1254 => x"5473802e",
  1255 => x"8a388c15",
  1256 => x"ff155555",
  1257 => x"a7990482",
  1258 => x"0bb0e40c",
  1259 => x"718f06b0",
  1260 => x"e00c81eb",
  1261 => x"51a3842d",
  1262 => x"b0d00881",
  1263 => x"2a708106",
  1264 => x"51527180",
  1265 => x"2ead3874",
  1266 => x"08852e09",
  1267 => x"8106a438",
  1268 => x"881580f5",
  1269 => x"2dff0552",
  1270 => x"71881681",
  1271 => x"b72d7198",
  1272 => x"2b527180",
  1273 => x"25883880",
  1274 => x"0b881681",
  1275 => x"b72d7451",
  1276 => x"a3e72d81",
  1277 => x"f451a384",
  1278 => x"2db0d008",
  1279 => x"812a7081",
  1280 => x"06515271",
  1281 => x"802eb338",
  1282 => x"7408852e",
  1283 => x"098106aa",
  1284 => x"38881580",
  1285 => x"f52d8105",
  1286 => x"52718816",
  1287 => x"81b72d71",
  1288 => x"81ff068b",
  1289 => x"1680f52d",
  1290 => x"54527272",
  1291 => x"27873872",
  1292 => x"881681b7",
  1293 => x"2d7451a3",
  1294 => x"e72d80da",
  1295 => x"51a3842d",
  1296 => x"b0d00881",
  1297 => x"2a708106",
  1298 => x"51527180",
  1299 => x"2e80ff38",
  1300 => x"b7b008b7",
  1301 => x"b8085553",
  1302 => x"73802e8a",
  1303 => x"388c13ff",
  1304 => x"155553a8",
  1305 => x"d8047208",
  1306 => x"5271822e",
  1307 => x"a6387182",
  1308 => x"26893871",
  1309 => x"812ea938",
  1310 => x"a9ce0471",
  1311 => x"832eb138",
  1312 => x"71842e09",
  1313 => x"810680c6",
  1314 => x"38881308",
  1315 => x"51a5b22d",
  1316 => x"a9ce04b7",
  1317 => x"b8085188",
  1318 => x"13085271",
  1319 => x"2da9ce04",
  1320 => x"810b8814",
  1321 => x"082bb7ac",
  1322 => x"0832b7ac",
  1323 => x"0ca9cb04",
  1324 => x"881380f5",
  1325 => x"2d81058b",
  1326 => x"1480f52d",
  1327 => x"53547174",
  1328 => x"24833880",
  1329 => x"54738814",
  1330 => x"81b72da4",
  1331 => x"972d8054",
  1332 => x"800bb0e4",
  1333 => x"0c738f06",
  1334 => x"b0e00ca0",
  1335 => x"5273b7b8",
  1336 => x"082e0981",
  1337 => x"069838b7",
  1338 => x"b408ff05",
  1339 => x"74327009",
  1340 => x"81057072",
  1341 => x"079f2a91",
  1342 => x"71315151",
  1343 => x"53537151",
  1344 => x"82ee2d81",
  1345 => x"14548e74",
  1346 => x"25c638b0",
  1347 => x"cc085271",
  1348 => x"b0d00c02",
  1349 => x"94050d04",
  1350 => x"00ffffff",
  1351 => x"ff00ffff",
  1352 => x"ffff00ff",
  1353 => x"ffffff00",
  1354 => x"52657365",
  1355 => x"74000000",
  1356 => x"53617665",
  1357 => x"20736574",
  1358 => x"74696e67",
  1359 => x"73000000",
  1360 => x"5363616e",
  1361 => x"6c696e65",
  1362 => x"73000000",
  1363 => x"4c6f6164",
  1364 => x"20524f4d",
  1365 => x"20100000",
  1366 => x"45786974",
  1367 => x"00000000",
  1368 => x"50432045",
  1369 => x"6e67696e",
  1370 => x"65206d6f",
  1371 => x"64650000",
  1372 => x"54757262",
  1373 => x"6f677261",
  1374 => x"66782031",
  1375 => x"36206d6f",
  1376 => x"64650000",
  1377 => x"56474120",
  1378 => x"2d203331",
  1379 => x"4b487a2c",
  1380 => x"20363048",
  1381 => x"7a000000",
  1382 => x"5456202d",
  1383 => x"20343830",
  1384 => x"692c2036",
  1385 => x"30487a00",
  1386 => x"4261636b",
  1387 => x"00000000",
  1388 => x"46504741",
  1389 => x"50434520",
  1390 => x"43464700",
  1391 => x"4c6f6164",
  1392 => x"696e6720",
  1393 => x"524f4d0a",
  1394 => x"00000000",
  1395 => x"52656164",
  1396 => x"20666169",
  1397 => x"6c65640a",
  1398 => x"00000000",
  1399 => x"4c6f6164",
  1400 => x"696e6720",
  1401 => x"00000000",
  1402 => x"496e6974",
  1403 => x"69616c69",
  1404 => x"7a696e67",
  1405 => x"20534420",
  1406 => x"63617264",
  1407 => x"0a000000",
  1408 => x"46696c65",
  1409 => x"73797374",
  1410 => x"656d2065",
  1411 => x"72726f72",
  1412 => x"0a000000",
  1413 => x"4d535833",
  1414 => x"42494f53",
  1415 => x"53595300",
  1416 => x"524f4d20",
  1417 => x"6c6f6164",
  1418 => x"696e6720",
  1419 => x"6661696c",
  1420 => x"65640a00",
  1421 => x"43617264",
  1422 => x"20696e69",
  1423 => x"74206661",
  1424 => x"696c6564",
  1425 => x"0a000000",
  1426 => x"4d425220",
  1427 => x"6661696c",
  1428 => x"0a000000",
  1429 => x"46415431",
  1430 => x"36202020",
  1431 => x"00000000",
  1432 => x"46415433",
  1433 => x"32202020",
  1434 => x"00000000",
  1435 => x"4e6f2070",
  1436 => x"61727469",
  1437 => x"74696f6e",
  1438 => x"20736967",
  1439 => x"0a000000",
  1440 => x"42616420",
  1441 => x"70617274",
  1442 => x"0a000000",
  1443 => x"53444843",
  1444 => x"20657272",
  1445 => x"6f72210a",
  1446 => x"00000000",
  1447 => x"53442069",
  1448 => x"6e69742e",
  1449 => x"2e2e0a00",
  1450 => x"53442063",
  1451 => x"61726420",
  1452 => x"72657365",
  1453 => x"74206661",
  1454 => x"696c6564",
  1455 => x"210a0000",
  1456 => x"57726974",
  1457 => x"65206661",
  1458 => x"696c6564",
  1459 => x"0a000000",
  1460 => x"16200000",
  1461 => x"14200000",
  1462 => x"15200000",
  1463 => x"00000002",
  1464 => x"00000002",
  1465 => x"00001528",
  1466 => x"000004d0",
  1467 => x"00000002",
  1468 => x"00001530",
  1469 => x"000003a4",
  1470 => x"00000003",
  1471 => x"00001748",
  1472 => x"00000002",
  1473 => x"00000001",
  1474 => x"00001540",
  1475 => x"00000001",
  1476 => x"00000003",
  1477 => x"00001740",
  1478 => x"00000002",
  1479 => x"00000002",
  1480 => x"0000154c",
  1481 => x"00000533",
  1482 => x"00000002",
  1483 => x"00001558",
  1484 => x"000011d4",
  1485 => x"00000000",
  1486 => x"00000000",
  1487 => x"00000000",
  1488 => x"00001560",
  1489 => x"00001570",
  1490 => x"00001584",
  1491 => x"00001598",
  1492 => x"00000002",
  1493 => x"0000187c",
  1494 => x"000004d4",
  1495 => x"00000002",
  1496 => x"0000188c",
  1497 => x"000004d4",
  1498 => x"00000002",
  1499 => x"0000189c",
  1500 => x"000004d4",
  1501 => x"00000002",
  1502 => x"000018ac",
  1503 => x"000004d4",
  1504 => x"00000002",
  1505 => x"000018bc",
  1506 => x"000004d4",
  1507 => x"00000002",
  1508 => x"000018cc",
  1509 => x"000004d4",
  1510 => x"00000002",
  1511 => x"000018dc",
  1512 => x"000004d4",
  1513 => x"00000002",
  1514 => x"000018ec",
  1515 => x"000004d4",
  1516 => x"00000002",
  1517 => x"000018fc",
  1518 => x"000004d4",
  1519 => x"00000002",
  1520 => x"0000190c",
  1521 => x"000004d4",
  1522 => x"00000002",
  1523 => x"0000191c",
  1524 => x"000004d4",
  1525 => x"00000002",
  1526 => x"0000192c",
  1527 => x"000004d4",
  1528 => x"00000002",
  1529 => x"0000193c",
  1530 => x"000004d4",
  1531 => x"00000004",
  1532 => x"000015a8",
  1533 => x"000016e0",
  1534 => x"00000000",
  1535 => x"00000000",
  1536 => x"00000000",
  1537 => x"00000000",
  1538 => x"00000000",
  1539 => x"00000000",
  1540 => x"00000000",
  1541 => x"00000000",
  1542 => x"00000000",
  1543 => x"00000000",
  1544 => x"00000000",
  1545 => x"00000000",
  1546 => x"00000000",
  1547 => x"00000000",
  1548 => x"00000000",
  1549 => x"00000000",
  1550 => x"00000000",
  1551 => x"00000000",
  1552 => x"00000000",
  1553 => x"00000000",
  1554 => x"00000000",
  1555 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

