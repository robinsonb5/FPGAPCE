-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb5",
     9 => x"d0080b0b",
    10 => x"0bb5d408",
    11 => x"0b0b0bb5",
    12 => x"d8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b5d80c0b",
    16 => x"0b0bb5d4",
    17 => x"0c0b0b0b",
    18 => x"b5d00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bafc4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b5d070bc",
    57 => x"c8278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8cdd0402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b5e00c9f",
    65 => x"0bb5e40c",
    66 => x"a0717081",
    67 => x"055334b5",
    68 => x"e408ff05",
    69 => x"b5e40cb5",
    70 => x"e4088025",
    71 => x"eb38b5e0",
    72 => x"08ff05b5",
    73 => x"e00cb5e0",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb5e0",
    94 => x"08258f38",
    95 => x"82b22db5",
    96 => x"e008ff05",
    97 => x"b5e00c82",
    98 => x"f404b5e0",
    99 => x"08b5e408",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b5e008",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b5",
   108 => x"e4088105",
   109 => x"b5e40cb5",
   110 => x"e408519f",
   111 => x"7125e238",
   112 => x"800bb5e4",
   113 => x"0cb5e008",
   114 => x"8105b5e0",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b5e40881",
   120 => x"05b5e40c",
   121 => x"b5e408a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b5e40cb5",
   125 => x"e0088105",
   126 => x"b5e00c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb5",
   155 => x"e80cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb5e8",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b5e80884",
   167 => x"07b5e80c",
   168 => x"5573842b",
   169 => x"87e87125",
   170 => x"83713170",
   171 => x"0b0b0bb2",
   172 => x"d80c8171",
   173 => x"2bf6880c",
   174 => x"fea413ff",
   175 => x"122c7888",
   176 => x"29ff9405",
   177 => x"70812cb5",
   178 => x"e8085258",
   179 => x"52555152",
   180 => x"5476802e",
   181 => x"85387081",
   182 => x"075170f6",
   183 => x"940c7109",
   184 => x"8105f680",
   185 => x"0c720981",
   186 => x"05f6840c",
   187 => x"0294050d",
   188 => x"0402f405",
   189 => x"0d745372",
   190 => x"70810554",
   191 => x"80f52d52",
   192 => x"71802e89",
   193 => x"38715182",
   194 => x"ee2d85f7",
   195 => x"04028c05",
   196 => x"0d0402f4",
   197 => x"050d7470",
   198 => x"8206bcb0",
   199 => x"0cb2f471",
   200 => x"81065454",
   201 => x"51718814",
   202 => x"81b72d70",
   203 => x"822a7081",
   204 => x"06515170",
   205 => x"941481b7",
   206 => x"2d70b5d0",
   207 => x"0c028c05",
   208 => x"0d0402f4",
   209 => x"050db0dc",
   210 => x"52b5f051",
   211 => x"95fb2db5",
   212 => x"d008802e",
   213 => x"9538b7d0",
   214 => x"52b5f051",
   215 => x"98b12db7",
   216 => x"d00870fe",
   217 => x"c00c5186",
   218 => x"922d028c",
   219 => x"050d0402",
   220 => x"f8050dbc",
   221 => x"b0088206",
   222 => x"b2fc0b80",
   223 => x"f52d5252",
   224 => x"70802e85",
   225 => x"38718107",
   226 => x"52b3940b",
   227 => x"80f52d51",
   228 => x"70802e85",
   229 => x"38718407",
   230 => x"52b5fc08",
   231 => x"802e8538",
   232 => x"71900752",
   233 => x"71b5d00c",
   234 => x"0288050d",
   235 => x"0402f005",
   236 => x"0d86ef2d",
   237 => x"b5d008b0",
   238 => x"dc53b5f0",
   239 => x"525395fb",
   240 => x"2db5d008",
   241 => x"802ea338",
   242 => x"72b7d00c",
   243 => x"b7d45480",
   244 => x"fd538074",
   245 => x"70840556",
   246 => x"0cff1353",
   247 => x"728025f2",
   248 => x"38b7d052",
   249 => x"b5f05198",
   250 => x"d72d0290",
   251 => x"050d0402",
   252 => x"d8050d81",
   253 => x"0bfec40c",
   254 => x"840bfec4",
   255 => x"0c7b52b5",
   256 => x"f05195fb",
   257 => x"2db5d008",
   258 => x"53b5d008",
   259 => x"802e81c7",
   260 => x"38b5f408",
   261 => x"56800bff",
   262 => x"17585976",
   263 => x"792e8b38",
   264 => x"81197781",
   265 => x"2a585976",
   266 => x"f738f719",
   267 => x"769fff06",
   268 => x"54597280",
   269 => x"2e8b38fc",
   270 => x"8016b5f0",
   271 => x"52569884",
   272 => x"2d75b080",
   273 => x"802e0981",
   274 => x"068f3886",
   275 => x"ef2db5d0",
   276 => x"088807fe",
   277 => x"c00c88e1",
   278 => x"04815380",
   279 => x"762580fd",
   280 => x"38785276",
   281 => x"5184802d",
   282 => x"b7d052b5",
   283 => x"f05198b1",
   284 => x"2db5d008",
   285 => x"b7d05b53",
   286 => x"8058b5d0",
   287 => x"08b03889",
   288 => x"c1047970",
   289 => x"84055b08",
   290 => x"7083fe80",
   291 => x"0671882b",
   292 => x"83fe8006",
   293 => x"71882a07",
   294 => x"72882a83",
   295 => x"fe800673",
   296 => x"982a07fe",
   297 => x"c80cfec8",
   298 => x"0c568419",
   299 => x"59537553",
   300 => x"84807625",
   301 => x"84388480",
   302 => x"53727824",
   303 => x"c53889c7",
   304 => x"04b0e851",
   305 => x"89da04b5",
   306 => x"f0519884",
   307 => x"2dfc8016",
   308 => x"81185856",
   309 => x"88d904b0",
   310 => x"f85185f1",
   311 => x"2d72b5d0",
   312 => x"0c02a805",
   313 => x"0d0402fc",
   314 => x"050da5c5",
   315 => x"2dfec451",
   316 => x"81710c82",
   317 => x"710c0284",
   318 => x"050d0402",
   319 => x"f4050d74",
   320 => x"10157084",
   321 => x"29b3d005",
   322 => x"70085551",
   323 => x"5272802e",
   324 => x"9b387280",
   325 => x"f52d5271",
   326 => x"802e9138",
   327 => x"b1805185",
   328 => x"f12d7251",
   329 => x"85f12d72",
   330 => x"5187ef2d",
   331 => x"b2dc51a7",
   332 => x"a32da5c5",
   333 => x"2d805184",
   334 => x"e52d028c",
   335 => x"050d0402",
   336 => x"e8050d80",
   337 => x"70565675",
   338 => x"b5800825",
   339 => x"af38bbdc",
   340 => x"08762ea8",
   341 => x"38745195",
   342 => x"a62db5d0",
   343 => x"08098105",
   344 => x"70b5d008",
   345 => x"079f2a77",
   346 => x"05811757",
   347 => x"575275b5",
   348 => x"80082588",
   349 => x"38bbdc08",
   350 => x"7526da38",
   351 => x"805674bb",
   352 => x"dc082780",
   353 => x"d0387451",
   354 => x"95a62d75",
   355 => x"842b52b5",
   356 => x"d008802e",
   357 => x"ae38b680",
   358 => x"128117b5",
   359 => x"d0085657",
   360 => x"528a5373",
   361 => x"70810555",
   362 => x"80f52d72",
   363 => x"70810554",
   364 => x"81b72dff",
   365 => x"13537280",
   366 => x"25e93880",
   367 => x"7281b72d",
   368 => x"8bcc04b5",
   369 => x"d008b680",
   370 => x"1381b72d",
   371 => x"8115558b",
   372 => x"7625ffaa",
   373 => x"38029805",
   374 => x"0d0402fc",
   375 => x"050d7251",
   376 => x"70fd2ead",
   377 => x"3870fd24",
   378 => x"8a3870fc",
   379 => x"2e80c438",
   380 => x"8cbb0470",
   381 => x"fe2eb138",
   382 => x"70ff2e09",
   383 => x"8106bc38",
   384 => x"b5800851",
   385 => x"70802eb3",
   386 => x"38ff11b5",
   387 => x"800c8cbb",
   388 => x"04b58008",
   389 => x"f00570b5",
   390 => x"800c5170",
   391 => x"80259c38",
   392 => x"800bb580",
   393 => x"0c8cbb04",
   394 => x"b5800881",
   395 => x"05b5800c",
   396 => x"8cbb04b5",
   397 => x"80089005",
   398 => x"b5800c8a",
   399 => x"bf2da688",
   400 => x"2d028405",
   401 => x"0d0402fc",
   402 => x"050d800b",
   403 => x"b5800c8a",
   404 => x"bf2db3cc",
   405 => x"51a7a32d",
   406 => x"0284050d",
   407 => x"0402f405",
   408 => x"0d810bb5",
   409 => x"fc0c9051",
   410 => x"86922d81",
   411 => x"0bfec40c",
   412 => x"900bfec0",
   413 => x"0c840bfe",
   414 => x"c40c830b",
   415 => x"fecc0ca3",
   416 => x"932da5a6",
   417 => x"2da2f82d",
   418 => x"a2f82d81",
   419 => x"f72d8151",
   420 => x"84e52da2",
   421 => x"f82da2f8",
   422 => x"2d815184",
   423 => x"e52db18c",
   424 => x"5185f12d",
   425 => x"84529d8a",
   426 => x"2d8f942d",
   427 => x"b5d00880",
   428 => x"2e8638fe",
   429 => x"528dc004",
   430 => x"ff125271",
   431 => x"8024e738",
   432 => x"71802e81",
   433 => x"813886c2",
   434 => x"2db1a451",
   435 => x"87ef2db5",
   436 => x"d008802e",
   437 => x"8f38b2dc",
   438 => x"51a7a32d",
   439 => x"805184e5",
   440 => x"2d8dee04",
   441 => x"b5d00851",
   442 => x"8cc62da5",
   443 => x"b22da3ab",
   444 => x"2da7b32d",
   445 => x"b5d008bc",
   446 => x"b408882b",
   447 => x"bcb80807",
   448 => x"fed80c53",
   449 => x"86ef2db5",
   450 => x"d008b5ec",
   451 => x"082ea238",
   452 => x"b5d008b5",
   453 => x"ec0cb5d0",
   454 => x"08fec00c",
   455 => x"84527251",
   456 => x"84e52da2",
   457 => x"f82da2f8",
   458 => x"2dff1252",
   459 => x"718025ee",
   460 => x"3872802e",
   461 => x"89388a0b",
   462 => x"fec40c8d",
   463 => x"ee04820b",
   464 => x"fec40c8d",
   465 => x"ee04b1b0",
   466 => x"5185f12d",
   467 => x"800bb5d0",
   468 => x"0c028c05",
   469 => x"0d0402e8",
   470 => x"050d7779",
   471 => x"7b585555",
   472 => x"80537276",
   473 => x"25a33874",
   474 => x"70810556",
   475 => x"80f52d74",
   476 => x"70810556",
   477 => x"80f52d52",
   478 => x"5271712e",
   479 => x"86388151",
   480 => x"8f8b0481",
   481 => x"13538ee2",
   482 => x"04805170",
   483 => x"b5d00c02",
   484 => x"98050d04",
   485 => x"02d8050d",
   486 => x"800bbbd8",
   487 => x"0cb7d052",
   488 => x"80519ff2",
   489 => x"2db5d008",
   490 => x"54b5d008",
   491 => x"8c38b1c4",
   492 => x"5185f12d",
   493 => x"735594af",
   494 => x"04805681",
   495 => x"0bbbfc0c",
   496 => x"8853b1d0",
   497 => x"52b88651",
   498 => x"8ed62db5",
   499 => x"d008762e",
   500 => x"09810687",
   501 => x"38b5d008",
   502 => x"bbfc0c88",
   503 => x"53b1dc52",
   504 => x"b8a2518e",
   505 => x"d62db5d0",
   506 => x"088738b5",
   507 => x"d008bbfc",
   508 => x"0cbbfc08",
   509 => x"802e80f6",
   510 => x"38bb960b",
   511 => x"80f52dbb",
   512 => x"970b80f5",
   513 => x"2d71982b",
   514 => x"71902b07",
   515 => x"bb980b80",
   516 => x"f52d7088",
   517 => x"2b7207bb",
   518 => x"990b80f5",
   519 => x"2d7107bb",
   520 => x"ce0b80f5",
   521 => x"2dbbcf0b",
   522 => x"80f52d71",
   523 => x"882b0753",
   524 => x"5f54525a",
   525 => x"56575573",
   526 => x"81abaa2e",
   527 => x"0981068d",
   528 => x"387551a1",
   529 => x"922db5d0",
   530 => x"085690da",
   531 => x"047382d4",
   532 => x"d52e8738",
   533 => x"b1e85191",
   534 => x"9b04b7d0",
   535 => x"5275519f",
   536 => x"f22db5d0",
   537 => x"0855b5d0",
   538 => x"08802e83",
   539 => x"c2388853",
   540 => x"b1dc52b8",
   541 => x"a2518ed6",
   542 => x"2db5d008",
   543 => x"8938810b",
   544 => x"bbd80c91",
   545 => x"a1048853",
   546 => x"b1d052b8",
   547 => x"86518ed6",
   548 => x"2db5d008",
   549 => x"802e8a38",
   550 => x"b1fc5185",
   551 => x"f12d91fb",
   552 => x"04bbce0b",
   553 => x"80f52d54",
   554 => x"7380d52e",
   555 => x"09810680",
   556 => x"ca38bbcf",
   557 => x"0b80f52d",
   558 => x"547381aa",
   559 => x"2e098106",
   560 => x"ba38800b",
   561 => x"b7d00b80",
   562 => x"f52d5654",
   563 => x"7481e92e",
   564 => x"83388154",
   565 => x"7481eb2e",
   566 => x"8c388055",
   567 => x"73752e09",
   568 => x"810682cb",
   569 => x"38b7db0b",
   570 => x"80f52d55",
   571 => x"748d38b7",
   572 => x"dc0b80f5",
   573 => x"2d547382",
   574 => x"2e863880",
   575 => x"5594af04",
   576 => x"b7dd0b80",
   577 => x"f52d70bb",
   578 => x"d00cff05",
   579 => x"bbd40cb7",
   580 => x"de0b80f5",
   581 => x"2db7df0b",
   582 => x"80f52d58",
   583 => x"76057782",
   584 => x"80290570",
   585 => x"bbe00cb7",
   586 => x"e00b80f5",
   587 => x"2d70bbf4",
   588 => x"0cbbd808",
   589 => x"59575876",
   590 => x"802e81a3",
   591 => x"388853b1",
   592 => x"dc52b8a2",
   593 => x"518ed62d",
   594 => x"b5d00881",
   595 => x"e238bbd0",
   596 => x"0870842b",
   597 => x"bbdc0c70",
   598 => x"bbf00cb7",
   599 => x"f50b80f5",
   600 => x"2db7f40b",
   601 => x"80f52d71",
   602 => x"82802905",
   603 => x"b7f60b80",
   604 => x"f52d7084",
   605 => x"80802912",
   606 => x"b7f70b80",
   607 => x"f52d7081",
   608 => x"800a2912",
   609 => x"70bbf80c",
   610 => x"bbf40871",
   611 => x"29bbe008",
   612 => x"0570bbe4",
   613 => x"0cb7fd0b",
   614 => x"80f52db7",
   615 => x"fc0b80f5",
   616 => x"2d718280",
   617 => x"2905b7fe",
   618 => x"0b80f52d",
   619 => x"70848080",
   620 => x"2912b7ff",
   621 => x"0b80f52d",
   622 => x"70982b81",
   623 => x"f00a0672",
   624 => x"0570bbe8",
   625 => x"0cfe117e",
   626 => x"297705bb",
   627 => x"ec0c5259",
   628 => x"5243545e",
   629 => x"51525952",
   630 => x"5d575957",
   631 => x"94ad04b7",
   632 => x"e20b80f5",
   633 => x"2db7e10b",
   634 => x"80f52d71",
   635 => x"82802905",
   636 => x"70bbdc0c",
   637 => x"70a02983",
   638 => x"ff057089",
   639 => x"2a70bbf0",
   640 => x"0cb7e70b",
   641 => x"80f52db7",
   642 => x"e60b80f5",
   643 => x"2d718280",
   644 => x"290570bb",
   645 => x"f80c7b71",
   646 => x"291e70bb",
   647 => x"ec0c7dbb",
   648 => x"e80c7305",
   649 => x"bbe40c55",
   650 => x"5e515155",
   651 => x"55815574",
   652 => x"b5d00c02",
   653 => x"a8050d04",
   654 => x"02ec050d",
   655 => x"7670872c",
   656 => x"7180ff06",
   657 => x"555654bb",
   658 => x"d8088a38",
   659 => x"73882c74",
   660 => x"81ff0654",
   661 => x"55b7d052",
   662 => x"bbe00815",
   663 => x"519ff22d",
   664 => x"b5d00854",
   665 => x"b5d00880",
   666 => x"2eb338bb",
   667 => x"d808802e",
   668 => x"98387284",
   669 => x"29b7d005",
   670 => x"70085253",
   671 => x"a1922db5",
   672 => x"d008f00a",
   673 => x"0653959b",
   674 => x"047210b7",
   675 => x"d0057080",
   676 => x"e02d5253",
   677 => x"a1c22db5",
   678 => x"d0085372",
   679 => x"5473b5d0",
   680 => x"0c029405",
   681 => x"0d0402ec",
   682 => x"050d7670",
   683 => x"842cbbec",
   684 => x"0805718f",
   685 => x"06525553",
   686 => x"728938b7",
   687 => x"d0527351",
   688 => x"9ff22d72",
   689 => x"a029b7d0",
   690 => x"05548074",
   691 => x"80f52d54",
   692 => x"5572752e",
   693 => x"83388155",
   694 => x"7281e52e",
   695 => x"93387480",
   696 => x"2e8e388b",
   697 => x"1480f52d",
   698 => x"98065372",
   699 => x"802e8338",
   700 => x"805473b5",
   701 => x"d00c0294",
   702 => x"050d0402",
   703 => x"cc050d7e",
   704 => x"605e5a80",
   705 => x"0bbbe808",
   706 => x"bbec0859",
   707 => x"5c568058",
   708 => x"bbdc0878",
   709 => x"2e81ae38",
   710 => x"778f06a0",
   711 => x"17575473",
   712 => x"8f38b7d0",
   713 => x"52765181",
   714 => x"17579ff2",
   715 => x"2db7d056",
   716 => x"807680f5",
   717 => x"2d565474",
   718 => x"742e8338",
   719 => x"81547481",
   720 => x"e52e80f6",
   721 => x"38817075",
   722 => x"06555c73",
   723 => x"802e80ea",
   724 => x"388b1680",
   725 => x"f52d9806",
   726 => x"597880de",
   727 => x"388b537c",
   728 => x"5275518e",
   729 => x"d62db5d0",
   730 => x"0880cf38",
   731 => x"9c160851",
   732 => x"a1922db5",
   733 => x"d008841b",
   734 => x"0c9a1680",
   735 => x"e02d51a1",
   736 => x"c22db5d0",
   737 => x"08b5d008",
   738 => x"881c0cb5",
   739 => x"d0085555",
   740 => x"bbd80880",
   741 => x"2e983894",
   742 => x"1680e02d",
   743 => x"51a1c22d",
   744 => x"b5d00890",
   745 => x"2b83fff0",
   746 => x"0a067016",
   747 => x"51547388",
   748 => x"1b0c787a",
   749 => x"0c7b5497",
   750 => x"fb048118",
   751 => x"58bbdc08",
   752 => x"7826fed4",
   753 => x"38bbd808",
   754 => x"802eae38",
   755 => x"7a5194b8",
   756 => x"2db5d008",
   757 => x"b5d00880",
   758 => x"fffffff8",
   759 => x"06555b73",
   760 => x"80ffffff",
   761 => x"f82e9238",
   762 => x"b5d008fe",
   763 => x"05bbd008",
   764 => x"29bbe408",
   765 => x"0557968e",
   766 => x"04805473",
   767 => x"b5d00c02",
   768 => x"b4050d04",
   769 => x"02f4050d",
   770 => x"74700881",
   771 => x"05710c70",
   772 => x"08bbd408",
   773 => x"06535371",
   774 => x"8e388813",
   775 => x"085194b8",
   776 => x"2db5d008",
   777 => x"88140c81",
   778 => x"0bb5d00c",
   779 => x"028c050d",
   780 => x"0402f005",
   781 => x"0d758811",
   782 => x"08fe05bb",
   783 => x"d00829bb",
   784 => x"e4081172",
   785 => x"08bbd408",
   786 => x"06057955",
   787 => x"5354549f",
   788 => x"f22d0290",
   789 => x"050d0402",
   790 => x"f0050d75",
   791 => x"881108fe",
   792 => x"05bbd008",
   793 => x"29bbe408",
   794 => x"117208bb",
   795 => x"d4080605",
   796 => x"79555354",
   797 => x"549eb22d",
   798 => x"0290050d",
   799 => x"0402f405",
   800 => x"0dd45281",
   801 => x"ff720c71",
   802 => x"085381ff",
   803 => x"720c7288",
   804 => x"2b83fe80",
   805 => x"06720870",
   806 => x"81ff0651",
   807 => x"525381ff",
   808 => x"720c7271",
   809 => x"07882b72",
   810 => x"087081ff",
   811 => x"06515253",
   812 => x"81ff720c",
   813 => x"72710788",
   814 => x"2b720870",
   815 => x"81ff0672",
   816 => x"07b5d00c",
   817 => x"5253028c",
   818 => x"050d0402",
   819 => x"f4050d74",
   820 => x"767181ff",
   821 => x"06d40c53",
   822 => x"53bc8008",
   823 => x"85387189",
   824 => x"2b527198",
   825 => x"2ad40c71",
   826 => x"902a7081",
   827 => x"ff06d40c",
   828 => x"5171882a",
   829 => x"7081ff06",
   830 => x"d40c5171",
   831 => x"81ff06d4",
   832 => x"0c72902a",
   833 => x"7081ff06",
   834 => x"d40c51d4",
   835 => x"087081ff",
   836 => x"06515182",
   837 => x"b8bf5270",
   838 => x"81ff2e09",
   839 => x"81069438",
   840 => x"81ff0bd4",
   841 => x"0cd40870",
   842 => x"81ff06ff",
   843 => x"14545151",
   844 => x"71e53870",
   845 => x"b5d00c02",
   846 => x"8c050d04",
   847 => x"02fc050d",
   848 => x"81c75181",
   849 => x"ff0bd40c",
   850 => x"ff115170",
   851 => x"8025f438",
   852 => x"0284050d",
   853 => x"0402f005",
   854 => x"0d9abc2d",
   855 => x"8fcf5380",
   856 => x"5287fc80",
   857 => x"f75199cb",
   858 => x"2db5d008",
   859 => x"54b5d008",
   860 => x"812e0981",
   861 => x"06a33881",
   862 => x"ff0bd40c",
   863 => x"820a5284",
   864 => x"9c80e951",
   865 => x"99cb2db5",
   866 => x"d0088b38",
   867 => x"81ff0bd4",
   868 => x"0c73539b",
   869 => x"9f049abc",
   870 => x"2dff1353",
   871 => x"72c13872",
   872 => x"b5d00c02",
   873 => x"90050d04",
   874 => x"02f4050d",
   875 => x"81ff0bd4",
   876 => x"0c935380",
   877 => x"5287fc80",
   878 => x"c15199cb",
   879 => x"2db5d008",
   880 => x"8b3881ff",
   881 => x"0bd40c81",
   882 => x"539bd504",
   883 => x"9abc2dff",
   884 => x"135372df",
   885 => x"3872b5d0",
   886 => x"0c028c05",
   887 => x"0d0402f0",
   888 => x"050d9abc",
   889 => x"2d83aa52",
   890 => x"849c80c8",
   891 => x"5199cb2d",
   892 => x"b5d00881",
   893 => x"2e098106",
   894 => x"923898fd",
   895 => x"2db5d008",
   896 => x"83ffff06",
   897 => x"537283aa",
   898 => x"2e97389b",
   899 => x"a82d9c9c",
   900 => x"0481549d",
   901 => x"8104b288",
   902 => x"5185f12d",
   903 => x"80549d81",
   904 => x"0481ff0b",
   905 => x"d40cb153",
   906 => x"9ad52db5",
   907 => x"d008802e",
   908 => x"80c03880",
   909 => x"5287fc80",
   910 => x"fa5199cb",
   911 => x"2db5d008",
   912 => x"b13881ff",
   913 => x"0bd40cd4",
   914 => x"085381ff",
   915 => x"0bd40c81",
   916 => x"ff0bd40c",
   917 => x"81ff0bd4",
   918 => x"0c81ff0b",
   919 => x"d40c7286",
   920 => x"2a708106",
   921 => x"b5d00856",
   922 => x"51537280",
   923 => x"2e93389c",
   924 => x"91047282",
   925 => x"2eff9f38",
   926 => x"ff135372",
   927 => x"ffaa3872",
   928 => x"5473b5d0",
   929 => x"0c029005",
   930 => x"0d0402f0",
   931 => x"050d810b",
   932 => x"bc800c84",
   933 => x"54d00870",
   934 => x"8f2a7081",
   935 => x"06515153",
   936 => x"72f33872",
   937 => x"d00c9abc",
   938 => x"2db29851",
   939 => x"85f12dd0",
   940 => x"08708f2a",
   941 => x"70810651",
   942 => x"515372f3",
   943 => x"38810bd0",
   944 => x"0cb15380",
   945 => x"5284d480",
   946 => x"c05199cb",
   947 => x"2db5d008",
   948 => x"812ea138",
   949 => x"72822e09",
   950 => x"81068c38",
   951 => x"b2a45185",
   952 => x"f12d8053",
   953 => x"9ea904ff",
   954 => x"135372d7",
   955 => x"38ff1454",
   956 => x"73ffa238",
   957 => x"9bde2db5",
   958 => x"d008bc80",
   959 => x"0cb5d008",
   960 => x"8b388152",
   961 => x"87fc80d0",
   962 => x"5199cb2d",
   963 => x"81ff0bd4",
   964 => x"0cd00870",
   965 => x"8f2a7081",
   966 => x"06515153",
   967 => x"72f33872",
   968 => x"d00c81ff",
   969 => x"0bd40c81",
   970 => x"5372b5d0",
   971 => x"0c029005",
   972 => x"0d0402e8",
   973 => x"050d7856",
   974 => x"81ff0bd4",
   975 => x"0cd00870",
   976 => x"8f2a7081",
   977 => x"06515153",
   978 => x"72f33882",
   979 => x"810bd00c",
   980 => x"81ff0bd4",
   981 => x"0c775287",
   982 => x"fc80d851",
   983 => x"99cb2db5",
   984 => x"d008802e",
   985 => x"8c38b2bc",
   986 => x"5185f12d",
   987 => x"81539fe9",
   988 => x"0481ff0b",
   989 => x"d40c81fe",
   990 => x"0bd40c80",
   991 => x"ff557570",
   992 => x"84055708",
   993 => x"70982ad4",
   994 => x"0c70902c",
   995 => x"7081ff06",
   996 => x"d40c5470",
   997 => x"882c7081",
   998 => x"ff06d40c",
   999 => x"547081ff",
  1000 => x"06d40c54",
  1001 => x"ff155574",
  1002 => x"8025d338",
  1003 => x"81ff0bd4",
  1004 => x"0c81ff0b",
  1005 => x"d40c81ff",
  1006 => x"0bd40c86",
  1007 => x"8da05481",
  1008 => x"ff0bd40c",
  1009 => x"d40881ff",
  1010 => x"06557487",
  1011 => x"38ff1454",
  1012 => x"73ed3881",
  1013 => x"ff0bd40c",
  1014 => x"d008708f",
  1015 => x"2a708106",
  1016 => x"51515372",
  1017 => x"f33872d0",
  1018 => x"0c72b5d0",
  1019 => x"0c029805",
  1020 => x"0d0402e8",
  1021 => x"050d7855",
  1022 => x"805681ff",
  1023 => x"0bd40cd0",
  1024 => x"08708f2a",
  1025 => x"70810651",
  1026 => x"515372f3",
  1027 => x"3882810b",
  1028 => x"d00c81ff",
  1029 => x"0bd40c77",
  1030 => x"5287fc80",
  1031 => x"d15199cb",
  1032 => x"2d80dbc6",
  1033 => x"df54b5d0",
  1034 => x"08802e8a",
  1035 => x"38b0e851",
  1036 => x"85f12da1",
  1037 => x"890481ff",
  1038 => x"0bd40cd4",
  1039 => x"087081ff",
  1040 => x"06515372",
  1041 => x"81fe2e09",
  1042 => x"81069d38",
  1043 => x"80ff5398",
  1044 => x"fd2db5d0",
  1045 => x"08757084",
  1046 => x"05570cff",
  1047 => x"13537280",
  1048 => x"25ed3881",
  1049 => x"56a0ee04",
  1050 => x"ff145473",
  1051 => x"c93881ff",
  1052 => x"0bd40c81",
  1053 => x"ff0bd40c",
  1054 => x"d008708f",
  1055 => x"2a708106",
  1056 => x"51515372",
  1057 => x"f33872d0",
  1058 => x"0c75b5d0",
  1059 => x"0c029805",
  1060 => x"0d0402f4",
  1061 => x"050d7470",
  1062 => x"882a83fe",
  1063 => x"80067072",
  1064 => x"982a0772",
  1065 => x"882b87fc",
  1066 => x"80800673",
  1067 => x"982b81f0",
  1068 => x"0a067173",
  1069 => x"0707b5d0",
  1070 => x"0c565153",
  1071 => x"51028c05",
  1072 => x"0d0402f8",
  1073 => x"050d028e",
  1074 => x"0580f52d",
  1075 => x"74882b07",
  1076 => x"7083ffff",
  1077 => x"06b5d00c",
  1078 => x"51028805",
  1079 => x"0d0402fc",
  1080 => x"050d7251",
  1081 => x"80710c80",
  1082 => x"0b84120c",
  1083 => x"0284050d",
  1084 => x"0402f005",
  1085 => x"0d757008",
  1086 => x"84120853",
  1087 => x"5353ff54",
  1088 => x"71712ea8",
  1089 => x"38a5ac2d",
  1090 => x"84130870",
  1091 => x"84291488",
  1092 => x"11700870",
  1093 => x"81ff0684",
  1094 => x"18088111",
  1095 => x"8706841a",
  1096 => x"0c535155",
  1097 => x"515151a5",
  1098 => x"a62d7154",
  1099 => x"73b5d00c",
  1100 => x"0290050d",
  1101 => x"0402f805",
  1102 => x"0da5ac2d",
  1103 => x"e008708b",
  1104 => x"2a708106",
  1105 => x"51525270",
  1106 => x"802e9d38",
  1107 => x"bc840870",
  1108 => x"8429bc8c",
  1109 => x"057381ff",
  1110 => x"06710c51",
  1111 => x"51bc8408",
  1112 => x"81118706",
  1113 => x"bc840c51",
  1114 => x"800bbcac",
  1115 => x"0ca59f2d",
  1116 => x"a5a62d02",
  1117 => x"88050d04",
  1118 => x"02fc050d",
  1119 => x"a5ac2d81",
  1120 => x"0bbcac0c",
  1121 => x"a5a62dbc",
  1122 => x"ac085170",
  1123 => x"fa380284",
  1124 => x"050d0402",
  1125 => x"fc050dbc",
  1126 => x"8451a1de",
  1127 => x"2da2b551",
  1128 => x"a59b2da4",
  1129 => x"c52d0284",
  1130 => x"050d0402",
  1131 => x"f4050da4",
  1132 => x"ad04b5d0",
  1133 => x"0881f02e",
  1134 => x"09810689",
  1135 => x"38810bb5",
  1136 => x"c40ca4ad",
  1137 => x"04b5d008",
  1138 => x"81e02e09",
  1139 => x"81068938",
  1140 => x"810bb5c8",
  1141 => x"0ca4ad04",
  1142 => x"b5d00852",
  1143 => x"b5c80880",
  1144 => x"2e8838b5",
  1145 => x"d0088180",
  1146 => x"05527184",
  1147 => x"2c728f06",
  1148 => x"5353b5c4",
  1149 => x"08802e99",
  1150 => x"38728429",
  1151 => x"b5840572",
  1152 => x"1381712b",
  1153 => x"70097308",
  1154 => x"06730c51",
  1155 => x"5353a4a3",
  1156 => x"04728429",
  1157 => x"b5840572",
  1158 => x"1383712b",
  1159 => x"72080772",
  1160 => x"0c535380",
  1161 => x"0bb5c80c",
  1162 => x"800bb5c4",
  1163 => x"0cbc8451",
  1164 => x"a1f12db5",
  1165 => x"d008ff24",
  1166 => x"fef83880",
  1167 => x"0bb5d00c",
  1168 => x"028c050d",
  1169 => x"0402f805",
  1170 => x"0db58452",
  1171 => x"8f518072",
  1172 => x"70840554",
  1173 => x"0cff1151",
  1174 => x"708025f2",
  1175 => x"38028805",
  1176 => x"0d0402f0",
  1177 => x"050d7551",
  1178 => x"a5ac2d70",
  1179 => x"822cfc06",
  1180 => x"b5841172",
  1181 => x"109e0671",
  1182 => x"0870722a",
  1183 => x"70830682",
  1184 => x"742b7009",
  1185 => x"7406760c",
  1186 => x"54515657",
  1187 => x"535153a5",
  1188 => x"a62d71b5",
  1189 => x"d00c0290",
  1190 => x"050d0471",
  1191 => x"980c04ff",
  1192 => x"b008b5d0",
  1193 => x"0c04810b",
  1194 => x"ffb00c04",
  1195 => x"800bffb0",
  1196 => x"0c0402fc",
  1197 => x"050d810b",
  1198 => x"b5cc0c81",
  1199 => x"5184e52d",
  1200 => x"0284050d",
  1201 => x"0402fc05",
  1202 => x"0d800bb5",
  1203 => x"cc0c8051",
  1204 => x"84e52d02",
  1205 => x"84050d04",
  1206 => x"02ec050d",
  1207 => x"76548052",
  1208 => x"870b8815",
  1209 => x"80f52d56",
  1210 => x"53747224",
  1211 => x"8338a053",
  1212 => x"725182ee",
  1213 => x"2d81128b",
  1214 => x"1580f52d",
  1215 => x"54527272",
  1216 => x"25de3802",
  1217 => x"94050d04",
  1218 => x"02f0050d",
  1219 => x"bcbc0854",
  1220 => x"81f72d80",
  1221 => x"0bbcc00c",
  1222 => x"7308802e",
  1223 => x"81803882",
  1224 => x"0bb5e40c",
  1225 => x"bcc0088f",
  1226 => x"06b5e00c",
  1227 => x"73085271",
  1228 => x"832e9638",
  1229 => x"71832689",
  1230 => x"3871812e",
  1231 => x"af38a789",
  1232 => x"0471852e",
  1233 => x"9f38a789",
  1234 => x"04881480",
  1235 => x"f52d8415",
  1236 => x"08b2cc53",
  1237 => x"545285f1",
  1238 => x"2d718429",
  1239 => x"13700852",
  1240 => x"52a78d04",
  1241 => x"7351a5d8",
  1242 => x"2da78904",
  1243 => x"bcb00888",
  1244 => x"15082c70",
  1245 => x"81065152",
  1246 => x"71802e87",
  1247 => x"38b2d051",
  1248 => x"a78604b2",
  1249 => x"d45185f1",
  1250 => x"2d841408",
  1251 => x"5185f12d",
  1252 => x"bcc00881",
  1253 => x"05bcc00c",
  1254 => x"8c1454a6",
  1255 => x"98040290",
  1256 => x"050d0471",
  1257 => x"bcbc0ca6",
  1258 => x"882dbcc0",
  1259 => x"08ff05bc",
  1260 => x"c40c0402",
  1261 => x"ec050dbc",
  1262 => x"bc085580",
  1263 => x"f851a4e2",
  1264 => x"2db5d008",
  1265 => x"812a7081",
  1266 => x"06515271",
  1267 => x"9b388751",
  1268 => x"a4e22db5",
  1269 => x"d008812a",
  1270 => x"70810651",
  1271 => x"5271802e",
  1272 => x"b138a7e8",
  1273 => x"04a3ab2d",
  1274 => x"8751a4e2",
  1275 => x"2db5d008",
  1276 => x"f438a7f8",
  1277 => x"04a3ab2d",
  1278 => x"80f851a4",
  1279 => x"e22db5d0",
  1280 => x"08f338b5",
  1281 => x"cc088132",
  1282 => x"70b5cc0c",
  1283 => x"70525284",
  1284 => x"e52d800b",
  1285 => x"bcb40c80",
  1286 => x"0bbcb80c",
  1287 => x"b5cc0882",
  1288 => x"dd3880da",
  1289 => x"51a4e22d",
  1290 => x"b5d00880",
  1291 => x"2e8a38bc",
  1292 => x"b4088180",
  1293 => x"07bcb40c",
  1294 => x"80d951a4",
  1295 => x"e22db5d0",
  1296 => x"08802e8a",
  1297 => x"38bcb408",
  1298 => x"80c007bc",
  1299 => x"b40c8194",
  1300 => x"51a4e22d",
  1301 => x"b5d00880",
  1302 => x"2e8938bc",
  1303 => x"b4089007",
  1304 => x"bcb40c81",
  1305 => x"9151a4e2",
  1306 => x"2db5d008",
  1307 => x"802e8938",
  1308 => x"bcb408a0",
  1309 => x"07bcb40c",
  1310 => x"81f551a4",
  1311 => x"e22db5d0",
  1312 => x"08802e89",
  1313 => x"38bcb408",
  1314 => x"8107bcb4",
  1315 => x"0c81f251",
  1316 => x"a4e22db5",
  1317 => x"d008802e",
  1318 => x"8938bcb4",
  1319 => x"088207bc",
  1320 => x"b40c81eb",
  1321 => x"51a4e22d",
  1322 => x"b5d00880",
  1323 => x"2e8938bc",
  1324 => x"b4088407",
  1325 => x"bcb40c81",
  1326 => x"f451a4e2",
  1327 => x"2db5d008",
  1328 => x"802e8938",
  1329 => x"bcb40888",
  1330 => x"07bcb40c",
  1331 => x"80d851a4",
  1332 => x"e22db5d0",
  1333 => x"08802e8a",
  1334 => x"38bcb808",
  1335 => x"818007bc",
  1336 => x"b80c9251",
  1337 => x"a4e22db5",
  1338 => x"d008802e",
  1339 => x"8a38bcb8",
  1340 => x"0880c007",
  1341 => x"bcb80c94",
  1342 => x"51a4e22d",
  1343 => x"b5d00880",
  1344 => x"2e8938bc",
  1345 => x"b8089007",
  1346 => x"bcb80c91",
  1347 => x"51a4e22d",
  1348 => x"b5d00880",
  1349 => x"2e8938bc",
  1350 => x"b808a007",
  1351 => x"bcb80c9d",
  1352 => x"51a4e22d",
  1353 => x"b5d00880",
  1354 => x"2e8938bc",
  1355 => x"b8088107",
  1356 => x"bcb80c9b",
  1357 => x"51a4e22d",
  1358 => x"b5d00880",
  1359 => x"2e8938bc",
  1360 => x"b8088207",
  1361 => x"bcb80c9c",
  1362 => x"51a4e22d",
  1363 => x"b5d00880",
  1364 => x"2e8938bc",
  1365 => x"b8088407",
  1366 => x"bcb80ca3",
  1367 => x"51a4e22d",
  1368 => x"b5d00880",
  1369 => x"2e8938bc",
  1370 => x"b8088807",
  1371 => x"bcb80c81",
  1372 => x"fd51a4e2",
  1373 => x"2d81fa51",
  1374 => x"a4e22daf",
  1375 => x"b90481f5",
  1376 => x"51a4e22d",
  1377 => x"b5d00881",
  1378 => x"2a708106",
  1379 => x"51527180",
  1380 => x"2eaf38bc",
  1381 => x"c4085271",
  1382 => x"802e8938",
  1383 => x"ff12bcc4",
  1384 => x"0cabc104",
  1385 => x"bcc00810",
  1386 => x"bcc00805",
  1387 => x"70842916",
  1388 => x"51528812",
  1389 => x"08802e89",
  1390 => x"38ff5188",
  1391 => x"12085271",
  1392 => x"2d81f251",
  1393 => x"a4e22db5",
  1394 => x"d008812a",
  1395 => x"70810651",
  1396 => x"5271802e",
  1397 => x"b138bcc0",
  1398 => x"08ff11bc",
  1399 => x"c4085653",
  1400 => x"53737225",
  1401 => x"89388114",
  1402 => x"bcc40cac",
  1403 => x"86047210",
  1404 => x"13708429",
  1405 => x"16515288",
  1406 => x"1208802e",
  1407 => x"8938fe51",
  1408 => x"88120852",
  1409 => x"712d81fd",
  1410 => x"51a4e22d",
  1411 => x"b5d00881",
  1412 => x"2a708106",
  1413 => x"51527180",
  1414 => x"2e863880",
  1415 => x"0bbcc40c",
  1416 => x"81fa51a4",
  1417 => x"e22db5d0",
  1418 => x"08812a70",
  1419 => x"81065152",
  1420 => x"71802e89",
  1421 => x"38bcc008",
  1422 => x"ff05bcc4",
  1423 => x"0cbcc408",
  1424 => x"70535473",
  1425 => x"802e8a38",
  1426 => x"8c15ff15",
  1427 => x"5555acc3",
  1428 => x"04820bb5",
  1429 => x"e40c718f",
  1430 => x"06b5e00c",
  1431 => x"81eb51a4",
  1432 => x"e22db5d0",
  1433 => x"08812a70",
  1434 => x"81065152",
  1435 => x"71802ead",
  1436 => x"38740885",
  1437 => x"2e098106",
  1438 => x"a4388815",
  1439 => x"80f52dff",
  1440 => x"05527188",
  1441 => x"1681b72d",
  1442 => x"71982b52",
  1443 => x"71802588",
  1444 => x"38800b88",
  1445 => x"1681b72d",
  1446 => x"7451a5d8",
  1447 => x"2d81f451",
  1448 => x"a4e22db5",
  1449 => x"d008812a",
  1450 => x"70810651",
  1451 => x"5271802e",
  1452 => x"b3387408",
  1453 => x"852e0981",
  1454 => x"06aa3888",
  1455 => x"1580f52d",
  1456 => x"81055271",
  1457 => x"881681b7",
  1458 => x"2d7181ff",
  1459 => x"068b1680",
  1460 => x"f52d5452",
  1461 => x"72722787",
  1462 => x"38728816",
  1463 => x"81b72d74",
  1464 => x"51a5d82d",
  1465 => x"80da51a4",
  1466 => x"e22db5d0",
  1467 => x"08812a70",
  1468 => x"81065152",
  1469 => x"71802e80",
  1470 => x"ff38bcbc",
  1471 => x"08bcc408",
  1472 => x"55537380",
  1473 => x"2e8a388c",
  1474 => x"13ff1555",
  1475 => x"53ae8204",
  1476 => x"72085271",
  1477 => x"822ea638",
  1478 => x"71822689",
  1479 => x"3871812e",
  1480 => x"a938aef8",
  1481 => x"0471832e",
  1482 => x"b1387184",
  1483 => x"2e098106",
  1484 => x"80c63888",
  1485 => x"130851a7",
  1486 => x"a32daef8",
  1487 => x"04bcc408",
  1488 => x"51881308",
  1489 => x"52712dae",
  1490 => x"f804810b",
  1491 => x"8814082b",
  1492 => x"bcb00832",
  1493 => x"bcb00cae",
  1494 => x"f5048813",
  1495 => x"80f52d81",
  1496 => x"058b1480",
  1497 => x"f52d5354",
  1498 => x"71742483",
  1499 => x"38805473",
  1500 => x"881481b7",
  1501 => x"2da6882d",
  1502 => x"8054800b",
  1503 => x"b5e40c73",
  1504 => x"8f06b5e0",
  1505 => x"0ca05273",
  1506 => x"bcc4082e",
  1507 => x"09810698",
  1508 => x"38bcc008",
  1509 => x"ff057432",
  1510 => x"70098105",
  1511 => x"7072079f",
  1512 => x"2a917131",
  1513 => x"51515353",
  1514 => x"715182ee",
  1515 => x"2d811454",
  1516 => x"8e7425c6",
  1517 => x"38b5cc08",
  1518 => x"5271b5d0",
  1519 => x"0c029405",
  1520 => x"0d040000",
  1521 => x"00ffffff",
  1522 => x"ff00ffff",
  1523 => x"ffff00ff",
  1524 => x"ffffff00",
  1525 => x"52657365",
  1526 => x"74000000",
  1527 => x"53617665",
  1528 => x"20736574",
  1529 => x"74696e67",
  1530 => x"73000000",
  1531 => x"5363616e",
  1532 => x"6c696e65",
  1533 => x"73000000",
  1534 => x"4c6f6164",
  1535 => x"20524f4d",
  1536 => x"20100000",
  1537 => x"45786974",
  1538 => x"00000000",
  1539 => x"50432045",
  1540 => x"6e67696e",
  1541 => x"65206d6f",
  1542 => x"64650000",
  1543 => x"54757262",
  1544 => x"6f677261",
  1545 => x"66782031",
  1546 => x"36206d6f",
  1547 => x"64650000",
  1548 => x"56474120",
  1549 => x"2d203331",
  1550 => x"4b487a2c",
  1551 => x"20363048",
  1552 => x"7a000000",
  1553 => x"5456202d",
  1554 => x"20343830",
  1555 => x"692c2036",
  1556 => x"30487a00",
  1557 => x"4261636b",
  1558 => x"00000000",
  1559 => x"46504741",
  1560 => x"50434520",
  1561 => x"43464700",
  1562 => x"52656164",
  1563 => x"20666169",
  1564 => x"6c65640a",
  1565 => x"00000000",
  1566 => x"4661696c",
  1567 => x"65640a00",
  1568 => x"4c6f6164",
  1569 => x"696e6720",
  1570 => x"00000000",
  1571 => x"496e6974",
  1572 => x"69616c69",
  1573 => x"7a696e67",
  1574 => x"20534420",
  1575 => x"63617264",
  1576 => x"0a000000",
  1577 => x"424f4f54",
  1578 => x"20202020",
  1579 => x"50434500",
  1580 => x"43617264",
  1581 => x"20696e69",
  1582 => x"74206661",
  1583 => x"696c6564",
  1584 => x"0a000000",
  1585 => x"4d425220",
  1586 => x"6661696c",
  1587 => x"0a000000",
  1588 => x"46415431",
  1589 => x"36202020",
  1590 => x"00000000",
  1591 => x"46415433",
  1592 => x"32202020",
  1593 => x"00000000",
  1594 => x"4e6f2070",
  1595 => x"61727469",
  1596 => x"74696f6e",
  1597 => x"20736967",
  1598 => x"0a000000",
  1599 => x"42616420",
  1600 => x"70617274",
  1601 => x"0a000000",
  1602 => x"53444843",
  1603 => x"20657272",
  1604 => x"6f72210a",
  1605 => x"00000000",
  1606 => x"53442069",
  1607 => x"6e69742e",
  1608 => x"2e2e0a00",
  1609 => x"53442063",
  1610 => x"61726420",
  1611 => x"72657365",
  1612 => x"74206661",
  1613 => x"696c6564",
  1614 => x"210a0000",
  1615 => x"57726974",
  1616 => x"65206661",
  1617 => x"696c6564",
  1618 => x"0a000000",
  1619 => x"16200000",
  1620 => x"14200000",
  1621 => x"15200000",
  1622 => x"00000002",
  1623 => x"00000002",
  1624 => x"000017d4",
  1625 => x"000004e6",
  1626 => x"00000002",
  1627 => x"000017dc",
  1628 => x"000003ad",
  1629 => x"00000003",
  1630 => x"000019c4",
  1631 => x"00000002",
  1632 => x"00000001",
  1633 => x"000017ec",
  1634 => x"00000002",
  1635 => x"00000003",
  1636 => x"000019bc",
  1637 => x"00000002",
  1638 => x"00000002",
  1639 => x"000017f8",
  1640 => x"00000646",
  1641 => x"00000002",
  1642 => x"00001804",
  1643 => x"000012c5",
  1644 => x"00000000",
  1645 => x"00000000",
  1646 => x"00000000",
  1647 => x"0000180c",
  1648 => x"0000181c",
  1649 => x"00001830",
  1650 => x"00001844",
  1651 => x"00000002",
  1652 => x"00001b00",
  1653 => x"000004fb",
  1654 => x"00000002",
  1655 => x"00001b10",
  1656 => x"000004fb",
  1657 => x"00000002",
  1658 => x"00001b20",
  1659 => x"000004fb",
  1660 => x"00000002",
  1661 => x"00001b30",
  1662 => x"000004fb",
  1663 => x"00000002",
  1664 => x"00001b40",
  1665 => x"000004fb",
  1666 => x"00000002",
  1667 => x"00001b50",
  1668 => x"000004fb",
  1669 => x"00000002",
  1670 => x"00001b60",
  1671 => x"000004fb",
  1672 => x"00000002",
  1673 => x"00001b70",
  1674 => x"000004fb",
  1675 => x"00000002",
  1676 => x"00001b80",
  1677 => x"000004fb",
  1678 => x"00000002",
  1679 => x"00001b90",
  1680 => x"000004fb",
  1681 => x"00000002",
  1682 => x"00001ba0",
  1683 => x"000004fb",
  1684 => x"00000002",
  1685 => x"00001bb0",
  1686 => x"000004fb",
  1687 => x"00000002",
  1688 => x"00001bc0",
  1689 => x"000004fb",
  1690 => x"00000004",
  1691 => x"00001854",
  1692 => x"0000195c",
  1693 => x"00000000",
  1694 => x"00000000",
  1695 => x"000005da",
  1696 => x"00000000",
  1697 => x"00000000",
  1698 => x"00000000",
  1699 => x"00000000",
  1700 => x"00000000",
  1701 => x"00000000",
  1702 => x"00000000",
  1703 => x"00000000",
  1704 => x"00000000",
  1705 => x"00000000",
  1706 => x"00000000",
  1707 => x"00000000",
  1708 => x"00000000",
  1709 => x"00000000",
  1710 => x"00000000",
  1711 => x"00000000",
  1712 => x"00000000",
  1713 => x"00000000",
  1714 => x"00000000",
  1715 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

