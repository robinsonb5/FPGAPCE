-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb7",
     9 => x"f8080b0b",
    10 => x"0bb7fc08",
    11 => x"0b0b0bb8",
    12 => x"80080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b8800c0b",
    16 => x"0b0bb7fc",
    17 => x"0c0b0b0b",
    18 => x"b7f80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0baed8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b7f870bd",
    57 => x"b0278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8d9a0402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b8880c9f",
    65 => x"0bb88c0c",
    66 => x"a0717081",
    67 => x"055334b8",
    68 => x"8c08ff05",
    69 => x"b88c0cb8",
    70 => x"8c088025",
    71 => x"eb38b888",
    72 => x"08ff05b8",
    73 => x"880cb888",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb888",
    94 => x"08258f38",
    95 => x"82b22db8",
    96 => x"8808ff05",
    97 => x"b8880c82",
    98 => x"f404b888",
    99 => x"08b88c08",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b88808",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b8",
   108 => x"8c088105",
   109 => x"b88c0cb8",
   110 => x"8c08519f",
   111 => x"7125e238",
   112 => x"800bb88c",
   113 => x"0cb88808",
   114 => x"8105b888",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b88c0881",
   120 => x"05b88c0c",
   121 => x"b88c08a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b88c0cb8",
   125 => x"88088105",
   126 => x"b8880c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb8",
   155 => x"900cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb890",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b8900884",
   167 => x"07b8900c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0bb4",
   172 => x"d80c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cb89008",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f8050d",
   198 => x"a68f2d80",
   199 => x"da51a7c6",
   200 => x"2db7f808",
   201 => x"812a7081",
   202 => x"06515271",
   203 => x"802ee938",
   204 => x"0288050d",
   205 => x"0402f405",
   206 => x"0dbda008",
   207 => x"99c406b6",
   208 => x"d40b80f5",
   209 => x"2d525270",
   210 => x"802e8638",
   211 => x"71848007",
   212 => x"52b68c0b",
   213 => x"80f52d72",
   214 => x"07b6b00b",
   215 => x"80f52d70",
   216 => x"812a7081",
   217 => x"06515354",
   218 => x"5270802e",
   219 => x"86387182",
   220 => x"80075272",
   221 => x"81065170",
   222 => x"802e8538",
   223 => x"71880752",
   224 => x"b6bc0b80",
   225 => x"f52d7084",
   226 => x"2b730781",
   227 => x"8432b7f8",
   228 => x"0c51028c",
   229 => x"050d0402",
   230 => x"f4050d74",
   231 => x"70818432",
   232 => x"bda00c70",
   233 => x"83065253",
   234 => x"70b6840b",
   235 => x"880581b7",
   236 => x"2d72892a",
   237 => x"70810651",
   238 => x"5170b6d4",
   239 => x"0b81b72d",
   240 => x"72832a81",
   241 => x"0673882a",
   242 => x"70810651",
   243 => x"52527080",
   244 => x"2e853871",
   245 => x"82075271",
   246 => x"b6b00b81",
   247 => x"b72d7284",
   248 => x"2c708306",
   249 => x"515170b6",
   250 => x"bc0b81b7",
   251 => x"2d70b7f8",
   252 => x"0c028c05",
   253 => x"0d0402f4",
   254 => x"050db5bc",
   255 => x"0b881180",
   256 => x"f52d8c12",
   257 => x"881180f5",
   258 => x"2d70842b",
   259 => x"73078c13",
   260 => x"881180f5",
   261 => x"2d70882b",
   262 => x"73079413",
   263 => x"80f52d70",
   264 => x"8c2b7207",
   265 => x"b7f80c53",
   266 => x"53535353",
   267 => x"56525351",
   268 => x"028c050d",
   269 => x"0402f405",
   270 => x"0d74b5bc",
   271 => x"71870655",
   272 => x"53517288",
   273 => x"1381b72d",
   274 => x"8c127184",
   275 => x"2c708706",
   276 => x"55525272",
   277 => x"881381b7",
   278 => x"2d8c1271",
   279 => x"842c7087",
   280 => x"06555252",
   281 => x"72881381",
   282 => x"b72d7084",
   283 => x"2c708706",
   284 => x"51517094",
   285 => x"1381b72d",
   286 => x"028c050d",
   287 => x"0402d405",
   288 => x"0d7cb1d8",
   289 => x"525585f3",
   290 => x"2d9dc02d",
   291 => x"b7f80880",
   292 => x"2e83ad38",
   293 => x"86b52db7",
   294 => x"f8085390",
   295 => x"892db7f8",
   296 => x"0854b7f8",
   297 => x"08802e83",
   298 => x"9938a1c3",
   299 => x"2db7f808",
   300 => x"802e8738",
   301 => x"b1f05189",
   302 => x"c70499ac",
   303 => x"2db7f808",
   304 => x"802ea238",
   305 => x"b2845185",
   306 => x"f32db29c",
   307 => x"5185f32d",
   308 => x"86942d72",
   309 => x"84075381",
   310 => x"0bfec40c",
   311 => x"72fec00c",
   312 => x"72518797",
   313 => x"2d840bfe",
   314 => x"c40cb2b8",
   315 => x"52b89851",
   316 => x"969b2db7",
   317 => x"f808802e",
   318 => x"80ec3874",
   319 => x"822e0981",
   320 => x"06af3872",
   321 => x"b8a40c87",
   322 => x"f62db7f8",
   323 => x"08b8a80c",
   324 => x"b8ac5480",
   325 => x"fd538074",
   326 => x"70840556",
   327 => x"0cff1353",
   328 => x"728025f2",
   329 => x"38b8a452",
   330 => x"b8985199",
   331 => x"862d8ae6",
   332 => x"0474812e",
   333 => x"098106ae",
   334 => x"38b2b852",
   335 => x"b8985196",
   336 => x"9b2db7f8",
   337 => x"08802e9e",
   338 => x"38b8a452",
   339 => x"b8985198",
   340 => x"e02db8a4",
   341 => x"08b8a808",
   342 => x"525388b5",
   343 => x"2d72fec0",
   344 => x"0c725187",
   345 => x"972db2c4",
   346 => x"5185f32d",
   347 => x"b2dc52b8",
   348 => x"9851969b",
   349 => x"2db7f808",
   350 => x"9838b2e8",
   351 => x"5185f32d",
   352 => x"b38052b8",
   353 => x"9851969b",
   354 => x"2db7f808",
   355 => x"802e81b0",
   356 => x"38b38c51",
   357 => x"85f32db8",
   358 => x"9c085780",
   359 => x"77595a76",
   360 => x"7a2e8b38",
   361 => x"811a7881",
   362 => x"2a595a77",
   363 => x"f738f71a",
   364 => x"5a807725",
   365 => x"81803879",
   366 => x"52775184",
   367 => x"802db8a4",
   368 => x"52b89851",
   369 => x"98e02db7",
   370 => x"f80853b7",
   371 => x"f808802e",
   372 => x"80c938b8",
   373 => x"a45b8059",
   374 => x"8c88047a",
   375 => x"7084055c",
   376 => x"087081ff",
   377 => x"0671882c",
   378 => x"7081ff06",
   379 => x"73902c70",
   380 => x"81ff0675",
   381 => x"982afec8",
   382 => x"0cfec80c",
   383 => x"58fec80c",
   384 => x"57fec80c",
   385 => x"841a5a53",
   386 => x"76538480",
   387 => x"77258438",
   388 => x"84805372",
   389 => x"7924c438",
   390 => x"8ca604b3",
   391 => x"9c5185f3",
   392 => x"2d72548c",
   393 => x"c204b898",
   394 => x"5198b32d",
   395 => x"fc801781",
   396 => x"1959578b",
   397 => x"b104820b",
   398 => x"fec40c81",
   399 => x"548cc204",
   400 => x"805473b7",
   401 => x"f80c02ac",
   402 => x"050d0402",
   403 => x"f8050da8",
   404 => x"962d81f7",
   405 => x"2d815184",
   406 => x"e52dfec4",
   407 => x"5281720c",
   408 => x"a58f2da5",
   409 => x"8f2d8472",
   410 => x"0c735188",
   411 => x"fd2db4dc",
   412 => x"51a9f42d",
   413 => x"805184e5",
   414 => x"2d028805",
   415 => x"0d0402fc",
   416 => x"050d8251",
   417 => x"8ccb2d02",
   418 => x"84050d04",
   419 => x"02fc050d",
   420 => x"80518ccb",
   421 => x"2d028405",
   422 => x"0d0402ec",
   423 => x"050d84b8",
   424 => x"5187972d",
   425 => x"810bfec4",
   426 => x"0c84b80b",
   427 => x"fec00c84",
   428 => x"0bfec40c",
   429 => x"830bfecc",
   430 => x"0ca5aa2d",
   431 => x"a88a2da5",
   432 => x"8f2da58f",
   433 => x"2d81f72d",
   434 => x"815184e5",
   435 => x"2da58f2d",
   436 => x"a58f2d81",
   437 => x"5184e52d",
   438 => x"815188fd",
   439 => x"2db7f808",
   440 => x"802e81d2",
   441 => x"38805184",
   442 => x"e52db4dc",
   443 => x"51a9f42d",
   444 => x"bd800889",
   445 => x"38bd8408",
   446 => x"802e80e2",
   447 => x"38fed008",
   448 => x"70810651",
   449 => x"5271802e",
   450 => x"80d438a8",
   451 => x"902dbd80",
   452 => x"0870bd84",
   453 => x"08705755",
   454 => x"565280ff",
   455 => x"72258438",
   456 => x"80ff5280",
   457 => x"ff732584",
   458 => x"3880ff53",
   459 => x"71ff8025",
   460 => x"8438ff80",
   461 => x"5272ff80",
   462 => x"258438ff",
   463 => x"80537472",
   464 => x"31bd800c",
   465 => x"737331bd",
   466 => x"840ca88a",
   467 => x"2d71882b",
   468 => x"83fe8006",
   469 => x"7381ff06",
   470 => x"7107fed0",
   471 => x"0c52a68f",
   472 => x"2daa842d",
   473 => x"b7f80853",
   474 => x"86b52db7",
   475 => x"f808fec0",
   476 => x"0c87f62d",
   477 => x"b7f808fe",
   478 => x"d40c86b5",
   479 => x"2db7f808",
   480 => x"b894082e",
   481 => x"9c38b7f8",
   482 => x"08b8940c",
   483 => x"84527251",
   484 => x"84e52da5",
   485 => x"8f2da58f",
   486 => x"2dff1252",
   487 => x"718025ee",
   488 => x"3872802e",
   489 => x"89388a0b",
   490 => x"fec40c8d",
   491 => x"f004820b",
   492 => x"fec40c8d",
   493 => x"f004b3ac",
   494 => x"5185f32d",
   495 => x"820bfec4",
   496 => x"0c800bb7",
   497 => x"f80c0294",
   498 => x"050d0402",
   499 => x"e8050d77",
   500 => x"797b5855",
   501 => x"55805372",
   502 => x"7625a338",
   503 => x"74708105",
   504 => x"5680f52d",
   505 => x"74708105",
   506 => x"5680f52d",
   507 => x"52527171",
   508 => x"2e863881",
   509 => x"51908004",
   510 => x"8113538f",
   511 => x"d7048051",
   512 => x"70b7f80c",
   513 => x"0298050d",
   514 => x"0402d805",
   515 => x"0d800bbc",
   516 => x"ac0cb8a4",
   517 => x"528051a0",
   518 => x"a82db7f8",
   519 => x"0854b7f8",
   520 => x"088c38b3",
   521 => x"c45185f3",
   522 => x"2d735595",
   523 => x"a4048056",
   524 => x"810bbcd0",
   525 => x"0c8853b3",
   526 => x"d052b8da",
   527 => x"518fcb2d",
   528 => x"b7f80876",
   529 => x"2e098106",
   530 => x"8738b7f8",
   531 => x"08bcd00c",
   532 => x"8853b3dc",
   533 => x"52b8f651",
   534 => x"8fcb2db7",
   535 => x"f8088738",
   536 => x"b7f808bc",
   537 => x"d00cbcd0",
   538 => x"08802e80",
   539 => x"f638bbea",
   540 => x"0b80f52d",
   541 => x"bbeb0b80",
   542 => x"f52d7198",
   543 => x"2b71902b",
   544 => x"07bbec0b",
   545 => x"80f52d70",
   546 => x"882b7207",
   547 => x"bbed0b80",
   548 => x"f52d7107",
   549 => x"bca20b80",
   550 => x"f52dbca3",
   551 => x"0b80f52d",
   552 => x"71882b07",
   553 => x"535f5452",
   554 => x"5a565755",
   555 => x"7381abaa",
   556 => x"2e098106",
   557 => x"8d387551",
   558 => x"a1ca2db7",
   559 => x"f8085691",
   560 => x"cf047382",
   561 => x"d4d52e87",
   562 => x"38b3e851",
   563 => x"929004b8",
   564 => x"a4527551",
   565 => x"a0a82db7",
   566 => x"f80855b7",
   567 => x"f808802e",
   568 => x"83c23888",
   569 => x"53b3dc52",
   570 => x"b8f6518f",
   571 => x"cb2db7f8",
   572 => x"08893881",
   573 => x"0bbcac0c",
   574 => x"92960488",
   575 => x"53b3d052",
   576 => x"b8da518f",
   577 => x"cb2db7f8",
   578 => x"08802e8a",
   579 => x"38b3fc51",
   580 => x"85f32d92",
   581 => x"f004bca2",
   582 => x"0b80f52d",
   583 => x"547380d5",
   584 => x"2e098106",
   585 => x"80ca38bc",
   586 => x"a30b80f5",
   587 => x"2d547381",
   588 => x"aa2e0981",
   589 => x"06ba3880",
   590 => x"0bb8a40b",
   591 => x"80f52d56",
   592 => x"547481e9",
   593 => x"2e833881",
   594 => x"547481eb",
   595 => x"2e8c3880",
   596 => x"5573752e",
   597 => x"09810682",
   598 => x"cb38b8af",
   599 => x"0b80f52d",
   600 => x"55748d38",
   601 => x"b8b00b80",
   602 => x"f52d5473",
   603 => x"822e8638",
   604 => x"805595a4",
   605 => x"04b8b10b",
   606 => x"80f52d70",
   607 => x"bca40cff",
   608 => x"05bca80c",
   609 => x"b8b20b80",
   610 => x"f52db8b3",
   611 => x"0b80f52d",
   612 => x"58760577",
   613 => x"82802905",
   614 => x"70bcb00c",
   615 => x"b8b40b80",
   616 => x"f52d70bc",
   617 => x"c40cbcac",
   618 => x"08595758",
   619 => x"76802e81",
   620 => x"a3388853",
   621 => x"b3dc52b8",
   622 => x"f6518fcb",
   623 => x"2db7f808",
   624 => x"81e238bc",
   625 => x"a4087084",
   626 => x"2bbcc80c",
   627 => x"70bcc00c",
   628 => x"b8c90b80",
   629 => x"f52db8c8",
   630 => x"0b80f52d",
   631 => x"71828029",
   632 => x"05b8ca0b",
   633 => x"80f52d70",
   634 => x"84808029",
   635 => x"12b8cb0b",
   636 => x"80f52d70",
   637 => x"81800a29",
   638 => x"1270bccc",
   639 => x"0cbcc408",
   640 => x"7129bcb0",
   641 => x"080570bc",
   642 => x"b40cb8d1",
   643 => x"0b80f52d",
   644 => x"b8d00b80",
   645 => x"f52d7182",
   646 => x"802905b8",
   647 => x"d20b80f5",
   648 => x"2d708480",
   649 => x"802912b8",
   650 => x"d30b80f5",
   651 => x"2d70982b",
   652 => x"81f00a06",
   653 => x"720570bc",
   654 => x"b80cfe11",
   655 => x"7e297705",
   656 => x"bcbc0c52",
   657 => x"59524354",
   658 => x"5e515259",
   659 => x"525d5759",
   660 => x"5795a204",
   661 => x"b8b60b80",
   662 => x"f52db8b5",
   663 => x"0b80f52d",
   664 => x"71828029",
   665 => x"0570bcc8",
   666 => x"0c70a029",
   667 => x"83ff0570",
   668 => x"892a70bc",
   669 => x"c00cb8bb",
   670 => x"0b80f52d",
   671 => x"b8ba0b80",
   672 => x"f52d7182",
   673 => x"80290570",
   674 => x"bccc0c7b",
   675 => x"71291e70",
   676 => x"bcbc0c7d",
   677 => x"bcb80c73",
   678 => x"05bcb40c",
   679 => x"555e5151",
   680 => x"55558155",
   681 => x"74b7f80c",
   682 => x"02a8050d",
   683 => x"0402ec05",
   684 => x"0d767087",
   685 => x"2c7180ff",
   686 => x"06555654",
   687 => x"bcac088a",
   688 => x"3873882c",
   689 => x"7481ff06",
   690 => x"5455b8a4",
   691 => x"52bcb008",
   692 => x"1551a0a8",
   693 => x"2db7f808",
   694 => x"54b7f808",
   695 => x"802eb338",
   696 => x"bcac0880",
   697 => x"2e983872",
   698 => x"8429b8a4",
   699 => x"05700852",
   700 => x"53a1ca2d",
   701 => x"b7f808f0",
   702 => x"0a065396",
   703 => x"90047210",
   704 => x"b8a40570",
   705 => x"80e02d52",
   706 => x"53a1fa2d",
   707 => x"b7f80853",
   708 => x"725473b7",
   709 => x"f80c0294",
   710 => x"050d0402",
   711 => x"c8050d7f",
   712 => x"615f5b80",
   713 => x"0bbcb808",
   714 => x"bcbc0859",
   715 => x"5d56bcac",
   716 => x"08762e8a",
   717 => x"38bca408",
   718 => x"842b5896",
   719 => x"c404bcc0",
   720 => x"08842b58",
   721 => x"80597878",
   722 => x"2781a938",
   723 => x"788f06a0",
   724 => x"17575473",
   725 => x"8f38b8a4",
   726 => x"52765181",
   727 => x"1757a0a8",
   728 => x"2db8a456",
   729 => x"807680f5",
   730 => x"2d565474",
   731 => x"742e8338",
   732 => x"81547481",
   733 => x"e52e80f6",
   734 => x"38817075",
   735 => x"06555d73",
   736 => x"802e80ea",
   737 => x"388b1680",
   738 => x"f52d9806",
   739 => x"5a7980de",
   740 => x"388b537d",
   741 => x"5275518f",
   742 => x"cb2db7f8",
   743 => x"0880cf38",
   744 => x"9c160851",
   745 => x"a1ca2db7",
   746 => x"f808841c",
   747 => x"0c9a1680",
   748 => x"e02d51a1",
   749 => x"fa2db7f8",
   750 => x"08b7f808",
   751 => x"881d0cb7",
   752 => x"f8085555",
   753 => x"bcac0880",
   754 => x"2e983894",
   755 => x"1680e02d",
   756 => x"51a1fa2d",
   757 => x"b7f80890",
   758 => x"2b83fff0",
   759 => x"0a067016",
   760 => x"51547388",
   761 => x"1c0c797b",
   762 => x"0c7c5498",
   763 => x"aa048119",
   764 => x"5996c604",
   765 => x"bcac0880",
   766 => x"2eae387b",
   767 => x"5195ad2d",
   768 => x"b7f808b7",
   769 => x"f80880ff",
   770 => x"fffff806",
   771 => x"555c7380",
   772 => x"fffffff8",
   773 => x"2e9238b7",
   774 => x"f808fe05",
   775 => x"bca40829",
   776 => x"bcb40805",
   777 => x"5796c404",
   778 => x"805473b7",
   779 => x"f80c02b8",
   780 => x"050d0402",
   781 => x"f4050d74",
   782 => x"70088105",
   783 => x"710c7008",
   784 => x"bca80806",
   785 => x"5353718e",
   786 => x"38881308",
   787 => x"5195ad2d",
   788 => x"b7f80888",
   789 => x"140c810b",
   790 => x"b7f80c02",
   791 => x"8c050d04",
   792 => x"02f0050d",
   793 => x"75881108",
   794 => x"fe05bca4",
   795 => x"0829bcb4",
   796 => x"08117208",
   797 => x"bca80806",
   798 => x"05795553",
   799 => x"5454a0a8",
   800 => x"2d029005",
   801 => x"0d0402f0",
   802 => x"050d7588",
   803 => x"1108fe05",
   804 => x"bca40829",
   805 => x"bcb40811",
   806 => x"7208bca8",
   807 => x"08060579",
   808 => x"55535454",
   809 => x"9ee82d02",
   810 => x"90050d04",
   811 => x"bcac08b7",
   812 => x"f80c0402",
   813 => x"f4050dd4",
   814 => x"5281ff72",
   815 => x"0c710853",
   816 => x"81ff720c",
   817 => x"72882b83",
   818 => x"fe800672",
   819 => x"087081ff",
   820 => x"06515253",
   821 => x"81ff720c",
   822 => x"72710788",
   823 => x"2b720870",
   824 => x"81ff0651",
   825 => x"525381ff",
   826 => x"720c7271",
   827 => x"07882b72",
   828 => x"087081ff",
   829 => x"067207b7",
   830 => x"f80c5253",
   831 => x"028c050d",
   832 => x"0402f405",
   833 => x"0d747671",
   834 => x"81ff06d4",
   835 => x"0c5353bc",
   836 => x"d4088538",
   837 => x"71892b52",
   838 => x"71982ad4",
   839 => x"0c71902a",
   840 => x"7081ff06",
   841 => x"d40c5171",
   842 => x"882a7081",
   843 => x"ff06d40c",
   844 => x"517181ff",
   845 => x"06d40c72",
   846 => x"902a7081",
   847 => x"ff06d40c",
   848 => x"51d40870",
   849 => x"81ff0651",
   850 => x"5182b8bf",
   851 => x"527081ff",
   852 => x"2e098106",
   853 => x"943881ff",
   854 => x"0bd40cd4",
   855 => x"087081ff",
   856 => x"06ff1454",
   857 => x"515171e5",
   858 => x"3870b7f8",
   859 => x"0c028c05",
   860 => x"0d0402fc",
   861 => x"050d81c7",
   862 => x"5181ff0b",
   863 => x"d40cff11",
   864 => x"51708025",
   865 => x"f4380284",
   866 => x"050d0402",
   867 => x"f0050d9a",
   868 => x"f22d8fcf",
   869 => x"53805287",
   870 => x"fc80f751",
   871 => x"9a812db7",
   872 => x"f80854b7",
   873 => x"f808812e",
   874 => x"098106a3",
   875 => x"3881ff0b",
   876 => x"d40c820a",
   877 => x"52849c80",
   878 => x"e9519a81",
   879 => x"2db7f808",
   880 => x"8b3881ff",
   881 => x"0bd40c73",
   882 => x"539bd504",
   883 => x"9af22dff",
   884 => x"135372c1",
   885 => x"3872b7f8",
   886 => x"0c029005",
   887 => x"0d0402f4",
   888 => x"050d81ff",
   889 => x"0bd40c93",
   890 => x"53805287",
   891 => x"fc80c151",
   892 => x"9a812db7",
   893 => x"f8088b38",
   894 => x"81ff0bd4",
   895 => x"0c81539c",
   896 => x"8b049af2",
   897 => x"2dff1353",
   898 => x"72df3872",
   899 => x"b7f80c02",
   900 => x"8c050d04",
   901 => x"02f0050d",
   902 => x"9af22d83",
   903 => x"aa52849c",
   904 => x"80c8519a",
   905 => x"812db7f8",
   906 => x"08812e09",
   907 => x"81069238",
   908 => x"99b32db7",
   909 => x"f80883ff",
   910 => x"ff065372",
   911 => x"83aa2e97",
   912 => x"389bde2d",
   913 => x"9cd20481",
   914 => x"549db704",
   915 => x"b4885185",
   916 => x"f32d8054",
   917 => x"9db70481",
   918 => x"ff0bd40c",
   919 => x"b1539b8b",
   920 => x"2db7f808",
   921 => x"802e80c0",
   922 => x"38805287",
   923 => x"fc80fa51",
   924 => x"9a812db7",
   925 => x"f808b138",
   926 => x"81ff0bd4",
   927 => x"0cd40853",
   928 => x"81ff0bd4",
   929 => x"0c81ff0b",
   930 => x"d40c81ff",
   931 => x"0bd40c81",
   932 => x"ff0bd40c",
   933 => x"72862a70",
   934 => x"8106b7f8",
   935 => x"08565153",
   936 => x"72802e93",
   937 => x"389cc704",
   938 => x"72822eff",
   939 => x"9f38ff13",
   940 => x"5372ffaa",
   941 => x"38725473",
   942 => x"b7f80c02",
   943 => x"90050d04",
   944 => x"02f0050d",
   945 => x"810bbcd4",
   946 => x"0c8454d0",
   947 => x"08708f2a",
   948 => x"70810651",
   949 => x"515372f3",
   950 => x"3872d00c",
   951 => x"9af22db4",
   952 => x"985185f3",
   953 => x"2dd00870",
   954 => x"8f2a7081",
   955 => x"06515153",
   956 => x"72f33881",
   957 => x"0bd00cb1",
   958 => x"53805284",
   959 => x"d480c051",
   960 => x"9a812db7",
   961 => x"f808812e",
   962 => x"a1387282",
   963 => x"2e098106",
   964 => x"8c38b4a4",
   965 => x"5185f32d",
   966 => x"80539edf",
   967 => x"04ff1353",
   968 => x"72d738ff",
   969 => x"145473ff",
   970 => x"a2389c94",
   971 => x"2db7f808",
   972 => x"bcd40cb7",
   973 => x"f8088b38",
   974 => x"815287fc",
   975 => x"80d0519a",
   976 => x"812d81ff",
   977 => x"0bd40cd0",
   978 => x"08708f2a",
   979 => x"70810651",
   980 => x"515372f3",
   981 => x"3872d00c",
   982 => x"81ff0bd4",
   983 => x"0c815372",
   984 => x"b7f80c02",
   985 => x"90050d04",
   986 => x"02e8050d",
   987 => x"785681ff",
   988 => x"0bd40cd0",
   989 => x"08708f2a",
   990 => x"70810651",
   991 => x"515372f3",
   992 => x"3882810b",
   993 => x"d00c81ff",
   994 => x"0bd40c77",
   995 => x"5287fc80",
   996 => x"d8519a81",
   997 => x"2db7f808",
   998 => x"802e8c38",
   999 => x"b4bc5185",
  1000 => x"f32d8153",
  1001 => x"a09f0481",
  1002 => x"ff0bd40c",
  1003 => x"81fe0bd4",
  1004 => x"0c80ff55",
  1005 => x"75708405",
  1006 => x"57087098",
  1007 => x"2ad40c70",
  1008 => x"902c7081",
  1009 => x"ff06d40c",
  1010 => x"5470882c",
  1011 => x"7081ff06",
  1012 => x"d40c5470",
  1013 => x"81ff06d4",
  1014 => x"0c54ff15",
  1015 => x"55748025",
  1016 => x"d33881ff",
  1017 => x"0bd40c81",
  1018 => x"ff0bd40c",
  1019 => x"81ff0bd4",
  1020 => x"0c868da0",
  1021 => x"5481ff0b",
  1022 => x"d40cd408",
  1023 => x"81ff0655",
  1024 => x"748738ff",
  1025 => x"145473ed",
  1026 => x"3881ff0b",
  1027 => x"d40cd008",
  1028 => x"708f2a70",
  1029 => x"81065151",
  1030 => x"5372f338",
  1031 => x"72d00c72",
  1032 => x"b7f80c02",
  1033 => x"98050d04",
  1034 => x"02e8050d",
  1035 => x"78558056",
  1036 => x"81ff0bd4",
  1037 => x"0cd00870",
  1038 => x"8f2a7081",
  1039 => x"06515153",
  1040 => x"72f33882",
  1041 => x"810bd00c",
  1042 => x"81ff0bd4",
  1043 => x"0c775287",
  1044 => x"fc80d151",
  1045 => x"9a812d80",
  1046 => x"dbc6df54",
  1047 => x"b7f80880",
  1048 => x"2e8a38b3",
  1049 => x"9c5185f3",
  1050 => x"2da1ba04",
  1051 => x"81ff0bd4",
  1052 => x"0cd40870",
  1053 => x"81ff0651",
  1054 => x"537281fe",
  1055 => x"2e098106",
  1056 => x"9d3880ff",
  1057 => x"5399b32d",
  1058 => x"b7f80875",
  1059 => x"70840557",
  1060 => x"0cff1353",
  1061 => x"728025ed",
  1062 => x"388156a1",
  1063 => x"a404ff14",
  1064 => x"5473c938",
  1065 => x"81ff0bd4",
  1066 => x"0cd00870",
  1067 => x"8f2a7081",
  1068 => x"06515153",
  1069 => x"72f33872",
  1070 => x"d00c75b7",
  1071 => x"f80c0298",
  1072 => x"050d04bc",
  1073 => x"d408b7f8",
  1074 => x"0c0402f4",
  1075 => x"050d7470",
  1076 => x"882a83fe",
  1077 => x"80067072",
  1078 => x"982a0772",
  1079 => x"882b87fc",
  1080 => x"80800673",
  1081 => x"982b81f0",
  1082 => x"0a067173",
  1083 => x"0707b7f8",
  1084 => x"0c565153",
  1085 => x"51028c05",
  1086 => x"0d0402f8",
  1087 => x"050d028e",
  1088 => x"0580f52d",
  1089 => x"74882b07",
  1090 => x"7083ffff",
  1091 => x"06b7f80c",
  1092 => x"51028805",
  1093 => x"0d0402fc",
  1094 => x"050d7251",
  1095 => x"80710c80",
  1096 => x"0b84120c",
  1097 => x"0284050d",
  1098 => x"0402f005",
  1099 => x"0d757008",
  1100 => x"84120853",
  1101 => x"5353ff54",
  1102 => x"71712ea8",
  1103 => x"38a8902d",
  1104 => x"84130870",
  1105 => x"84291488",
  1106 => x"11700870",
  1107 => x"81ff0684",
  1108 => x"18088111",
  1109 => x"8706841a",
  1110 => x"0c535155",
  1111 => x"515151a8",
  1112 => x"8a2d7154",
  1113 => x"73b7f80c",
  1114 => x"0290050d",
  1115 => x"0402f405",
  1116 => x"0da8902d",
  1117 => x"e008e408",
  1118 => x"718b2a70",
  1119 => x"81065153",
  1120 => x"54527080",
  1121 => x"2e9d38bc",
  1122 => x"d8087084",
  1123 => x"29bce005",
  1124 => x"7381ff06",
  1125 => x"710c5151",
  1126 => x"bcd80881",
  1127 => x"118706bc",
  1128 => x"d80c5172",
  1129 => x"8b2a7081",
  1130 => x"06515170",
  1131 => x"802e8192",
  1132 => x"38b7a808",
  1133 => x"8429bd8c",
  1134 => x"057381ff",
  1135 => x"06710c51",
  1136 => x"b7a80881",
  1137 => x"05b7a80c",
  1138 => x"850bb7a4",
  1139 => x"0cb7a808",
  1140 => x"b7a0082e",
  1141 => x"09810681",
  1142 => x"a638800b",
  1143 => x"b7a80cbd",
  1144 => x"9c08819b",
  1145 => x"38bd8c08",
  1146 => x"70097083",
  1147 => x"06fecc0c",
  1148 => x"5270852a",
  1149 => x"708106bd",
  1150 => x"84085551",
  1151 => x"52537080",
  1152 => x"2e8e38bd",
  1153 => x"9408fe80",
  1154 => x"3212bd84",
  1155 => x"0ca49704",
  1156 => x"bd940812",
  1157 => x"bd840c72",
  1158 => x"842a7081",
  1159 => x"06bd8008",
  1160 => x"54515170",
  1161 => x"802e9038",
  1162 => x"bd900881",
  1163 => x"ff321281",
  1164 => x"05bd800c",
  1165 => x"a4ff0471",
  1166 => x"bd900831",
  1167 => x"bd800ca4",
  1168 => x"ff04b7a4",
  1169 => x"08ff05b7",
  1170 => x"a40cb7a4",
  1171 => x"08ff2e09",
  1172 => x"8106ac38",
  1173 => x"b7a80880",
  1174 => x"2e923881",
  1175 => x"0bbd9c0c",
  1176 => x"870bb7a0",
  1177 => x"0831b7a0",
  1178 => x"0ca4fa04",
  1179 => x"bd9c0851",
  1180 => x"70802e86",
  1181 => x"38ff11bd",
  1182 => x"9c0c800b",
  1183 => x"b7a80c80",
  1184 => x"0bbd880c",
  1185 => x"a8832da8",
  1186 => x"8a2d028c",
  1187 => x"050d0402",
  1188 => x"fc050da8",
  1189 => x"902d810b",
  1190 => x"bd880ca8",
  1191 => x"8a2dbd88",
  1192 => x"085170fa",
  1193 => x"38028405",
  1194 => x"0d0402f8",
  1195 => x"050dbcd8",
  1196 => x"51a2962d",
  1197 => x"800bbd9c",
  1198 => x"0c830bb7",
  1199 => x"a00ce408",
  1200 => x"708c2a70",
  1201 => x"81065151",
  1202 => x"5271802e",
  1203 => x"8638840b",
  1204 => x"b7a00ce4",
  1205 => x"08708d2a",
  1206 => x"70810651",
  1207 => x"51527180",
  1208 => x"2e9f3887",
  1209 => x"0bb7a008",
  1210 => x"31b7a00c",
  1211 => x"e408708a",
  1212 => x"2a708106",
  1213 => x"51515271",
  1214 => x"802ef138",
  1215 => x"81f40be4",
  1216 => x"0ca2ed51",
  1217 => x"a7ff2da7",
  1218 => x"a92d0288",
  1219 => x"050d0402",
  1220 => x"f4050da7",
  1221 => x"9104b7f8",
  1222 => x"0881f02e",
  1223 => x"09810689",
  1224 => x"38810bb7",
  1225 => x"ec0ca791",
  1226 => x"04b7f808",
  1227 => x"81e02e09",
  1228 => x"81068938",
  1229 => x"810bb7f0",
  1230 => x"0ca79104",
  1231 => x"b7f80852",
  1232 => x"b7f00880",
  1233 => x"2e8838b7",
  1234 => x"f8088180",
  1235 => x"05527184",
  1236 => x"2c728f06",
  1237 => x"5353b7ec",
  1238 => x"08802e99",
  1239 => x"38728429",
  1240 => x"b7ac0572",
  1241 => x"1381712b",
  1242 => x"70097308",
  1243 => x"06730c51",
  1244 => x"5353a787",
  1245 => x"04728429",
  1246 => x"b7ac0572",
  1247 => x"1383712b",
  1248 => x"72080772",
  1249 => x"0c535380",
  1250 => x"0bb7f00c",
  1251 => x"800bb7ec",
  1252 => x"0cbcd851",
  1253 => x"a2a92db7",
  1254 => x"f808ff24",
  1255 => x"fef83880",
  1256 => x"0bb7f80c",
  1257 => x"028c050d",
  1258 => x"0402f805",
  1259 => x"0db7ac52",
  1260 => x"8f518072",
  1261 => x"70840554",
  1262 => x"0cff1151",
  1263 => x"708025f2",
  1264 => x"38028805",
  1265 => x"0d0402f0",
  1266 => x"050d7551",
  1267 => x"a8902d70",
  1268 => x"822cfc06",
  1269 => x"b7ac1172",
  1270 => x"109e0671",
  1271 => x"0870722a",
  1272 => x"70830682",
  1273 => x"742b7009",
  1274 => x"7406760c",
  1275 => x"54515657",
  1276 => x"535153a8",
  1277 => x"8a2d71b7",
  1278 => x"f80c0290",
  1279 => x"050d0471",
  1280 => x"980c04ff",
  1281 => x"b008b7f8",
  1282 => x"0c04810b",
  1283 => x"ffb00c04",
  1284 => x"800bffb0",
  1285 => x"0c0402fc",
  1286 => x"050d800b",
  1287 => x"b7f40c80",
  1288 => x"5184e52d",
  1289 => x"0284050d",
  1290 => x"0402ec05",
  1291 => x"0d765480",
  1292 => x"52870b88",
  1293 => x"1580f52d",
  1294 => x"56537472",
  1295 => x"248338a0",
  1296 => x"53725182",
  1297 => x"ee2d8112",
  1298 => x"8b1580f5",
  1299 => x"2d545272",
  1300 => x"7225de38",
  1301 => x"0294050d",
  1302 => x"0402f005",
  1303 => x"0dbda408",
  1304 => x"5481f72d",
  1305 => x"800bbda8",
  1306 => x"0c730880",
  1307 => x"2e818038",
  1308 => x"820bb88c",
  1309 => x"0cbda808",
  1310 => x"8f06b888",
  1311 => x"0c730852",
  1312 => x"71832e96",
  1313 => x"38718326",
  1314 => x"89387181",
  1315 => x"2eaf38a9",
  1316 => x"da047185",
  1317 => x"2e9f38a9",
  1318 => x"da048814",
  1319 => x"80f52d84",
  1320 => x"1508b4cc",
  1321 => x"53545285",
  1322 => x"f32d7184",
  1323 => x"29137008",
  1324 => x"5252a9de",
  1325 => x"047351a8",
  1326 => x"a92da9da",
  1327 => x"04bda008",
  1328 => x"8815082c",
  1329 => x"70810651",
  1330 => x"5271802e",
  1331 => x"8738b4d0",
  1332 => x"51a9d704",
  1333 => x"b4d45185",
  1334 => x"f32d8414",
  1335 => x"085185f3",
  1336 => x"2dbda808",
  1337 => x"8105bda8",
  1338 => x"0c8c1454",
  1339 => x"a8e90402",
  1340 => x"90050d04",
  1341 => x"71bda40c",
  1342 => x"a8d92dbd",
  1343 => x"a808ff05",
  1344 => x"bdac0c04",
  1345 => x"02ec050d",
  1346 => x"bda40855",
  1347 => x"80f851a7",
  1348 => x"c62db7f8",
  1349 => x"08812a70",
  1350 => x"81065152",
  1351 => x"719b3887",
  1352 => x"51a7c62d",
  1353 => x"b7f80881",
  1354 => x"2a708106",
  1355 => x"51527180",
  1356 => x"2eb138aa",
  1357 => x"b904a68f",
  1358 => x"2d8751a7",
  1359 => x"c62db7f8",
  1360 => x"08f438aa",
  1361 => x"c904a68f",
  1362 => x"2d80f851",
  1363 => x"a7c62db7",
  1364 => x"f808f338",
  1365 => x"b7f40881",
  1366 => x"3270b7f4",
  1367 => x"0c705252",
  1368 => x"84e52db7",
  1369 => x"f408a238",
  1370 => x"80da51a7",
  1371 => x"c62d81f5",
  1372 => x"51a7c62d",
  1373 => x"81f251a7",
  1374 => x"c62d81eb",
  1375 => x"51a7c62d",
  1376 => x"81f451a7",
  1377 => x"c62daecd",
  1378 => x"0481f551",
  1379 => x"a7c62db7",
  1380 => x"f808812a",
  1381 => x"70810651",
  1382 => x"5271802e",
  1383 => x"8f38bdac",
  1384 => x"08527180",
  1385 => x"2e8638ff",
  1386 => x"12bdac0c",
  1387 => x"81f251a7",
  1388 => x"c62db7f8",
  1389 => x"08812a70",
  1390 => x"81065152",
  1391 => x"71802e95",
  1392 => x"38bda808",
  1393 => x"ff05bdac",
  1394 => x"08545272",
  1395 => x"72258638",
  1396 => x"8113bdac",
  1397 => x"0cbdac08",
  1398 => x"70535473",
  1399 => x"802e8a38",
  1400 => x"8c15ff15",
  1401 => x"5555abdb",
  1402 => x"04820bb8",
  1403 => x"8c0c718f",
  1404 => x"06b8880c",
  1405 => x"81eb51a7",
  1406 => x"c62db7f8",
  1407 => x"08812a70",
  1408 => x"81065152",
  1409 => x"71802ead",
  1410 => x"38740885",
  1411 => x"2e098106",
  1412 => x"a4388815",
  1413 => x"80f52dff",
  1414 => x"05527188",
  1415 => x"1681b72d",
  1416 => x"71982b52",
  1417 => x"71802588",
  1418 => x"38800b88",
  1419 => x"1681b72d",
  1420 => x"7451a8a9",
  1421 => x"2d81f451",
  1422 => x"a7c62db7",
  1423 => x"f808812a",
  1424 => x"70810651",
  1425 => x"5271802e",
  1426 => x"b3387408",
  1427 => x"852e0981",
  1428 => x"06aa3888",
  1429 => x"1580f52d",
  1430 => x"81055271",
  1431 => x"881681b7",
  1432 => x"2d7181ff",
  1433 => x"068b1680",
  1434 => x"f52d5452",
  1435 => x"72722787",
  1436 => x"38728816",
  1437 => x"81b72d74",
  1438 => x"51a8a92d",
  1439 => x"80da51a7",
  1440 => x"c62db7f8",
  1441 => x"08812a70",
  1442 => x"81065152",
  1443 => x"71802e80",
  1444 => x"fb38bda4",
  1445 => x"08bdac08",
  1446 => x"55537380",
  1447 => x"2e8a388c",
  1448 => x"13ff1555",
  1449 => x"53ad9a04",
  1450 => x"72085271",
  1451 => x"822ea638",
  1452 => x"71822689",
  1453 => x"3871812e",
  1454 => x"a538ae8c",
  1455 => x"0471832e",
  1456 => x"ad387184",
  1457 => x"2e098106",
  1458 => x"80c23888",
  1459 => x"130851a9",
  1460 => x"f42dae8c",
  1461 => x"04881308",
  1462 => x"52712dae",
  1463 => x"8c04810b",
  1464 => x"8814082b",
  1465 => x"bda00832",
  1466 => x"bda00cae",
  1467 => x"89048813",
  1468 => x"80f52d81",
  1469 => x"058b1480",
  1470 => x"f52d5354",
  1471 => x"71742483",
  1472 => x"38805473",
  1473 => x"881481b7",
  1474 => x"2da8d92d",
  1475 => x"8054800b",
  1476 => x"b88c0c73",
  1477 => x"8f06b888",
  1478 => x"0ca05273",
  1479 => x"bdac082e",
  1480 => x"09810698",
  1481 => x"38bda808",
  1482 => x"ff057432",
  1483 => x"70098105",
  1484 => x"7072079f",
  1485 => x"2a917131",
  1486 => x"51515353",
  1487 => x"715182ee",
  1488 => x"2d811454",
  1489 => x"8e7425c6",
  1490 => x"38b7f408",
  1491 => x"5271b7f8",
  1492 => x"0c029405",
  1493 => x"0d040000",
  1494 => x"00ffffff",
  1495 => x"ff00ffff",
  1496 => x"ffff00ff",
  1497 => x"ffffff00",
  1498 => x"52657365",
  1499 => x"74000000",
  1500 => x"53617665",
  1501 => x"20616e64",
  1502 => x"20526573",
  1503 => x"65740000",
  1504 => x"4f707469",
  1505 => x"6f6e7320",
  1506 => x"10000000",
  1507 => x"536f756e",
  1508 => x"64201000",
  1509 => x"54757262",
  1510 => x"6f000000",
  1511 => x"4d6f7573",
  1512 => x"6520656d",
  1513 => x"756c6174",
  1514 => x"696f6e00",
  1515 => x"45786974",
  1516 => x"00000000",
  1517 => x"4d617374",
  1518 => x"65720000",
  1519 => x"4f504c4c",
  1520 => x"00000000",
  1521 => x"53434300",
  1522 => x"50534700",
  1523 => x"4261636b",
  1524 => x"00000000",
  1525 => x"5363616e",
  1526 => x"6c696e65",
  1527 => x"73000000",
  1528 => x"53442043",
  1529 => x"61726400",
  1530 => x"4a617061",
  1531 => x"6e657365",
  1532 => x"206b6579",
  1533 => x"206c6179",
  1534 => x"6f757400",
  1535 => x"32303438",
  1536 => x"4b422052",
  1537 => x"414d0000",
  1538 => x"34303936",
  1539 => x"4b422052",
  1540 => x"414d0000",
  1541 => x"536c323a",
  1542 => x"204e6f6e",
  1543 => x"65000000",
  1544 => x"536c323a",
  1545 => x"20455345",
  1546 => x"2d534343",
  1547 => x"20314d42",
  1548 => x"2f534343",
  1549 => x"2d490000",
  1550 => x"536c323a",
  1551 => x"20455345",
  1552 => x"2d52414d",
  1553 => x"20314d42",
  1554 => x"2f415343",
  1555 => x"49493800",
  1556 => x"536c323a",
  1557 => x"20455345",
  1558 => x"2d52414d",
  1559 => x"20314d42",
  1560 => x"2f415343",
  1561 => x"49493136",
  1562 => x"00000000",
  1563 => x"536c313a",
  1564 => x"204e6f6e",
  1565 => x"65000000",
  1566 => x"536c313a",
  1567 => x"20455345",
  1568 => x"2d534343",
  1569 => x"20314d42",
  1570 => x"2f534343",
  1571 => x"2d490000",
  1572 => x"536c313a",
  1573 => x"204d6567",
  1574 => x"6152414d",
  1575 => x"00000000",
  1576 => x"56474120",
  1577 => x"2d203331",
  1578 => x"4b487a2c",
  1579 => x"20363048",
  1580 => x"7a000000",
  1581 => x"56474120",
  1582 => x"2d203331",
  1583 => x"4b487a2c",
  1584 => x"20353048",
  1585 => x"7a000000",
  1586 => x"5456202d",
  1587 => x"20343830",
  1588 => x"692c2036",
  1589 => x"30487a00",
  1590 => x"496e6974",
  1591 => x"69616c69",
  1592 => x"7a696e67",
  1593 => x"20534420",
  1594 => x"63617264",
  1595 => x"0a000000",
  1596 => x"53444843",
  1597 => x"206e6f74",
  1598 => x"20737570",
  1599 => x"706f7274",
  1600 => x"65643b00",
  1601 => x"46617433",
  1602 => x"32206e6f",
  1603 => x"74207375",
  1604 => x"70706f72",
  1605 => x"7465643b",
  1606 => x"00000000",
  1607 => x"0a646973",
  1608 => x"61626c69",
  1609 => x"6e672053",
  1610 => x"44206361",
  1611 => x"72640a10",
  1612 => x"204f4b0a",
  1613 => x"00000000",
  1614 => x"4f434d53",
  1615 => x"58202020",
  1616 => x"43464700",
  1617 => x"54727969",
  1618 => x"6e67204d",
  1619 => x"53583342",
  1620 => x"494f532e",
  1621 => x"5359530a",
  1622 => x"00000000",
  1623 => x"4d535833",
  1624 => x"42494f53",
  1625 => x"53595300",
  1626 => x"54727969",
  1627 => x"6e672042",
  1628 => x"494f535f",
  1629 => x"4d32502e",
  1630 => x"524f4d0a",
  1631 => x"00000000",
  1632 => x"42494f53",
  1633 => x"5f4d3250",
  1634 => x"524f4d00",
  1635 => x"4c6f6164",
  1636 => x"696e6720",
  1637 => x"42494f53",
  1638 => x"0a000000",
  1639 => x"52656164",
  1640 => x"20666169",
  1641 => x"6c65640a",
  1642 => x"00000000",
  1643 => x"4c6f6164",
  1644 => x"696e6720",
  1645 => x"42494f53",
  1646 => x"20666169",
  1647 => x"6c65640a",
  1648 => x"00000000",
  1649 => x"4d425220",
  1650 => x"6661696c",
  1651 => x"0a000000",
  1652 => x"46415431",
  1653 => x"36202020",
  1654 => x"00000000",
  1655 => x"46415433",
  1656 => x"32202020",
  1657 => x"00000000",
  1658 => x"4e6f2070",
  1659 => x"61727469",
  1660 => x"74696f6e",
  1661 => x"20736967",
  1662 => x"0a000000",
  1663 => x"42616420",
  1664 => x"70617274",
  1665 => x"0a000000",
  1666 => x"53444843",
  1667 => x"20657272",
  1668 => x"6f72210a",
  1669 => x"00000000",
  1670 => x"53442069",
  1671 => x"6e69742e",
  1672 => x"2e2e0a00",
  1673 => x"53442063",
  1674 => x"61726420",
  1675 => x"72657365",
  1676 => x"74206661",
  1677 => x"696c6564",
  1678 => x"210a0000",
  1679 => x"57726974",
  1680 => x"65206661",
  1681 => x"696c6564",
  1682 => x"0a000000",
  1683 => x"16200000",
  1684 => x"14200000",
  1685 => x"15200000",
  1686 => x"00000002",
  1687 => x"00000002",
  1688 => x"00001768",
  1689 => x"0000068c",
  1690 => x"00000002",
  1691 => x"00001770",
  1692 => x"0000067e",
  1693 => x"00000004",
  1694 => x"00001780",
  1695 => x"00001b04",
  1696 => x"00000004",
  1697 => x"0000178c",
  1698 => x"00001abc",
  1699 => x"00000001",
  1700 => x"00001794",
  1701 => x"00000007",
  1702 => x"00000001",
  1703 => x"0000179c",
  1704 => x"0000000a",
  1705 => x"00000002",
  1706 => x"000017ac",
  1707 => x"00001416",
  1708 => x"00000000",
  1709 => x"00000000",
  1710 => x"00000000",
  1711 => x"00000005",
  1712 => x"000017b4",
  1713 => x"00000007",
  1714 => x"00000005",
  1715 => x"000017bc",
  1716 => x"00000007",
  1717 => x"00000005",
  1718 => x"000017c4",
  1719 => x"00000007",
  1720 => x"00000005",
  1721 => x"000017c8",
  1722 => x"00000007",
  1723 => x"00000004",
  1724 => x"000017cc",
  1725 => x"00001a5c",
  1726 => x"00000000",
  1727 => x"00000000",
  1728 => x"00000000",
  1729 => x"00000003",
  1730 => x"00001b94",
  1731 => x"00000003",
  1732 => x"00000001",
  1733 => x"000017d4",
  1734 => x"0000000b",
  1735 => x"00000001",
  1736 => x"000017e0",
  1737 => x"00000002",
  1738 => x"00000003",
  1739 => x"00001b88",
  1740 => x"00000003",
  1741 => x"00000003",
  1742 => x"00001b78",
  1743 => x"00000004",
  1744 => x"00000001",
  1745 => x"000017e8",
  1746 => x"00000006",
  1747 => x"00000003",
  1748 => x"00001b70",
  1749 => x"00000002",
  1750 => x"00000004",
  1751 => x"000017cc",
  1752 => x"00001a5c",
  1753 => x"00000000",
  1754 => x"00000000",
  1755 => x"00000000",
  1756 => x"000017fc",
  1757 => x"00001808",
  1758 => x"00001814",
  1759 => x"00001820",
  1760 => x"00001838",
  1761 => x"00001850",
  1762 => x"0000186c",
  1763 => x"00001878",
  1764 => x"00001890",
  1765 => x"000018a0",
  1766 => x"000018b4",
  1767 => x"000018c8",
  1768 => x"00000003",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"00000000",
  1786 => x"00000000",
  1787 => x"00000000",
  1788 => x"00000000",
  1789 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

