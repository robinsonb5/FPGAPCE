-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bba",
     9 => x"b0080b0b",
    10 => x"0bbab408",
    11 => x"0b0b0bba",
    12 => x"b8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bab80c0b",
    16 => x"0b0bbab4",
    17 => x"0c0b0b0b",
    18 => x"bab00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb4a0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bab07080",
    57 => x"c2ec278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"518f8e04",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbac00c",
    65 => x"9f0bbac4",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"bac408ff",
    69 => x"05bac40c",
    70 => x"bac40880",
    71 => x"25eb38ba",
    72 => x"c008ff05",
    73 => x"bac00cba",
    74 => x"c0088025",
    75 => x"d7380284",
    76 => x"050d0402",
    77 => x"f0050df8",
    78 => x"8053f8a0",
    79 => x"5483bf52",
    80 => x"73708105",
    81 => x"55335170",
    82 => x"73708105",
    83 => x"5534ff12",
    84 => x"52718025",
    85 => x"eb38fbc0",
    86 => x"539f52a0",
    87 => x"73708105",
    88 => x"5534ff12",
    89 => x"52718025",
    90 => x"f2380290",
    91 => x"050d0402",
    92 => x"f4050d74",
    93 => x"538e0bba",
    94 => x"c008258f",
    95 => x"3882b32d",
    96 => x"bac008ff",
    97 => x"05bac00c",
    98 => x"82f504ba",
    99 => x"c008bac4",
   100 => x"08535172",
   101 => x"8a2e0981",
   102 => x"06b73871",
   103 => x"51719f24",
   104 => x"a038bac0",
   105 => x"08a02911",
   106 => x"f8801151",
   107 => x"51a07134",
   108 => x"bac40881",
   109 => x"05bac40c",
   110 => x"bac40851",
   111 => x"9f7125e2",
   112 => x"38800bba",
   113 => x"c40cbac0",
   114 => x"088105ba",
   115 => x"c00c83e5",
   116 => x"0470a029",
   117 => x"12f88011",
   118 => x"51517271",
   119 => x"34bac408",
   120 => x"8105bac4",
   121 => x"0cbac408",
   122 => x"a02e0981",
   123 => x"068e3880",
   124 => x"0bbac40c",
   125 => x"bac00881",
   126 => x"05bac00c",
   127 => x"028c050d",
   128 => x"0402e805",
   129 => x"0d777956",
   130 => x"56880bfc",
   131 => x"1677712c",
   132 => x"8f065452",
   133 => x"54805372",
   134 => x"72259538",
   135 => x"7153fbe0",
   136 => x"14518771",
   137 => x"348114ff",
   138 => x"14545472",
   139 => x"f1387153",
   140 => x"f9157671",
   141 => x"2c870653",
   142 => x"5171802e",
   143 => x"8b38fbe0",
   144 => x"14517171",
   145 => x"34811454",
   146 => x"728e2495",
   147 => x"388f7331",
   148 => x"53fbe014",
   149 => x"51a07134",
   150 => x"8114ff14",
   151 => x"545472f1",
   152 => x"38029805",
   153 => x"0d0402ec",
   154 => x"050d800b",
   155 => x"bac80cf6",
   156 => x"8c08f690",
   157 => x"0871882c",
   158 => x"565481ff",
   159 => x"06527372",
   160 => x"25883871",
   161 => x"54820bba",
   162 => x"c80c7288",
   163 => x"2c7381ff",
   164 => x"06545574",
   165 => x"73258b38",
   166 => x"72bac808",
   167 => x"8407bac8",
   168 => x"0c557384",
   169 => x"2b87e871",
   170 => x"25837131",
   171 => x"700b0b0b",
   172 => x"b7a00c81",
   173 => x"712bf688",
   174 => x"0cfea413",
   175 => x"ff122c78",
   176 => x"8829ff94",
   177 => x"0570812c",
   178 => x"bac80852",
   179 => x"58525551",
   180 => x"52547680",
   181 => x"2e853870",
   182 => x"81075170",
   183 => x"f6940c71",
   184 => x"098105f6",
   185 => x"800c7209",
   186 => x"8105f684",
   187 => x"0c029405",
   188 => x"0d0402f4",
   189 => x"050d7453",
   190 => x"72708105",
   191 => x"5480f52d",
   192 => x"5271802e",
   193 => x"89387151",
   194 => x"82ef2d85",
   195 => x"f804028c",
   196 => x"050d0402",
   197 => x"f4050d74",
   198 => x"70820680",
   199 => x"c2d00cb7",
   200 => x"bc718106",
   201 => x"54545171",
   202 => x"881481b7",
   203 => x"2d70822a",
   204 => x"70810651",
   205 => x"5170a014",
   206 => x"81b72d70",
   207 => x"bab00c02",
   208 => x"8c050d04",
   209 => x"02f8050d",
   210 => x"b5b852ba",
   211 => x"cc5199c0",
   212 => x"2dbab008",
   213 => x"802e9d38",
   214 => x"bde852ba",
   215 => x"cc519bff",
   216 => x"2dbde808",
   217 => x"bad80cbd",
   218 => x"e808fec0",
   219 => x"0cbde808",
   220 => x"5186932d",
   221 => x"0288050d",
   222 => x"0402f005",
   223 => x"0db5b852",
   224 => x"bacc5199",
   225 => x"c02dbab0",
   226 => x"08802ea5",
   227 => x"38bad808",
   228 => x"bde80cbd",
   229 => x"ec5480fd",
   230 => x"53807470",
   231 => x"8405560c",
   232 => x"ff135372",
   233 => x"8025f238",
   234 => x"bde852ba",
   235 => x"cc519ca8",
   236 => x"2d029005",
   237 => x"0d0402d4",
   238 => x"050dbad8",
   239 => x"08fec00c",
   240 => x"810bfec4",
   241 => x"0c840bfe",
   242 => x"c40c7c52",
   243 => x"bacc5199",
   244 => x"c02dbab0",
   245 => x"0853bab0",
   246 => x"08802e81",
   247 => x"cc38bad0",
   248 => x"0856800b",
   249 => x"ff175859",
   250 => x"76792e8b",
   251 => x"38811977",
   252 => x"812a5859",
   253 => x"76f738f7",
   254 => x"19769fff",
   255 => x"06545972",
   256 => x"802e8b38",
   257 => x"fc8016ba",
   258 => x"cc52569b",
   259 => x"d12d75b0",
   260 => x"80802e09",
   261 => x"81068938",
   262 => x"820bfedc",
   263 => x"0c88b704",
   264 => x"75988080",
   265 => x"2e098106",
   266 => x"8938810b",
   267 => x"fedc0c88",
   268 => x"b704800b",
   269 => x"fedc0c81",
   270 => x"5b807625",
   271 => x"80e93878",
   272 => x"52765184",
   273 => x"812dbde8",
   274 => x"52bacc51",
   275 => x"9bff2dba",
   276 => x"b008802e",
   277 => x"bb38bde8",
   278 => x"5a83fc58",
   279 => x"79708405",
   280 => x"5b087083",
   281 => x"fe800671",
   282 => x"882b83fe",
   283 => x"80067188",
   284 => x"2a077288",
   285 => x"2a83fe80",
   286 => x"0673982a",
   287 => x"07fec80c",
   288 => x"fec80c56",
   289 => x"fc195953",
   290 => x"778025d0",
   291 => x"38899704",
   292 => x"bab0085b",
   293 => x"848056ba",
   294 => x"cc519bd1",
   295 => x"2dfc8016",
   296 => x"81185856",
   297 => x"88b9047a",
   298 => x"5372bab0",
   299 => x"0c02ac05",
   300 => x"0d0402fc",
   301 => x"050da9ad",
   302 => x"2dfec451",
   303 => x"81710c82",
   304 => x"710c0284",
   305 => x"050d0402",
   306 => x"f4050d74",
   307 => x"10157084",
   308 => x"29b8b005",
   309 => x"70085551",
   310 => x"5272802e",
   311 => x"90387280",
   312 => x"f52d5271",
   313 => x"802e8638",
   314 => x"725187b6",
   315 => x"2db7a451",
   316 => x"ab912da9",
   317 => x"ad2d8051",
   318 => x"84e62d02",
   319 => x"8c050d04",
   320 => x"02f4050d",
   321 => x"74765451",
   322 => x"8a527270",
   323 => x"81055480",
   324 => x"f52d7170",
   325 => x"81055381",
   326 => x"b72dff12",
   327 => x"52718025",
   328 => x"e9388071",
   329 => x"81b72d02",
   330 => x"8c050d04",
   331 => x"02e0050d",
   332 => x"80705557",
   333 => x"76b9e008",
   334 => x"25b13880",
   335 => x"c1f40877",
   336 => x"2ea93876",
   337 => x"5198e22d",
   338 => x"bab00809",
   339 => x"810570ba",
   340 => x"b008079f",
   341 => x"2a750581",
   342 => x"19595553",
   343 => x"73b9e008",
   344 => x"25893880",
   345 => x"c1f40877",
   346 => x"26d93880",
   347 => x"547680c1",
   348 => x"f4082781",
   349 => x"98387651",
   350 => x"98e22dba",
   351 => x"b008802e",
   352 => x"80ef38ba",
   353 => x"b0088b05",
   354 => x"80f52d70",
   355 => x"842a7081",
   356 => x"06811777",
   357 => x"1078842b",
   358 => x"5b545b51",
   359 => x"54557280",
   360 => x"2eaf3873",
   361 => x"15822b8c",
   362 => x"920bb8b4",
   363 => x"120c5375",
   364 => x"743110ba",
   365 => x"e0115454",
   366 => x"90737081",
   367 => x"055581b7",
   368 => x"2da07381",
   369 => x"b72dbab0",
   370 => x"0852bae2",
   371 => x"14518be9",
   372 => x"04731582",
   373 => x"2b89c70b",
   374 => x"b8b4120c",
   375 => x"53bab008",
   376 => x"52757431",
   377 => x"10bae005",
   378 => x"5177548a",
   379 => x"802d8c84",
   380 => x"04739029",
   381 => x"74317010",
   382 => x"bae00551",
   383 => x"53bab008",
   384 => x"7381b72d",
   385 => x"8117578b",
   386 => x"7425fee1",
   387 => x"3802a005",
   388 => x"0d0402e8",
   389 => x"050d7756",
   390 => x"8070b9e0",
   391 => x"08185456",
   392 => x"53727224",
   393 => x"b83880c1",
   394 => x"f408732e",
   395 => x"b0387251",
   396 => x"98e22dba",
   397 => x"b008bab0",
   398 => x"08098105",
   399 => x"70bab008",
   400 => x"079f2a77",
   401 => x"058116b9",
   402 => x"e0081a53",
   403 => x"56575354",
   404 => x"74722489",
   405 => x"3880c1f4",
   406 => x"087326d2",
   407 => x"389a1480",
   408 => x"e02d51a5",
   409 => x"a12dbab0",
   410 => x"08539cd1",
   411 => x"2dbab008",
   412 => x"802e9738",
   413 => x"941480e0",
   414 => x"2d51a5a1",
   415 => x"2dbab008",
   416 => x"902b83ff",
   417 => x"f00a0673",
   418 => x"07537251",
   419 => x"91c72d8a",
   420 => x"ac2da9f0",
   421 => x"2d029805",
   422 => x"0d0402fc",
   423 => x"050d7251",
   424 => x"70fd2ead",
   425 => x"3870fd24",
   426 => x"8a3870fc",
   427 => x"2e80c438",
   428 => x"8dfb0470",
   429 => x"fe2eb138",
   430 => x"70ff2e09",
   431 => x"8106bc38",
   432 => x"b9e00851",
   433 => x"70802eb3",
   434 => x"38ff11b9",
   435 => x"e00c8dfb",
   436 => x"04b9e008",
   437 => x"f00570b9",
   438 => x"e00c5170",
   439 => x"80259c38",
   440 => x"800bb9e0",
   441 => x"0c8dfb04",
   442 => x"b9e00881",
   443 => x"05b9e00c",
   444 => x"8dfb04b9",
   445 => x"e0089005",
   446 => x"b9e00c8a",
   447 => x"ac2da9f0",
   448 => x"2d028405",
   449 => x"0d0402fc",
   450 => x"050dbad8",
   451 => x"08fb06ba",
   452 => x"d80c7251",
   453 => x"89c72d02",
   454 => x"84050d04",
   455 => x"02fc050d",
   456 => x"bad80884",
   457 => x"07bad80c",
   458 => x"725189c7",
   459 => x"2d028405",
   460 => x"0d0402fc",
   461 => x"050d800b",
   462 => x"b9e00c8a",
   463 => x"ac2db8ac",
   464 => x"51ab912d",
   465 => x"b89451ab",
   466 => x"a42d0284",
   467 => x"050d0402",
   468 => x"f8050d80",
   469 => x"c2d00882",
   470 => x"06b7c40b",
   471 => x"80f52d52",
   472 => x"5270802e",
   473 => x"85387181",
   474 => x"0752b7dc",
   475 => x"0b80f52d",
   476 => x"5170802e",
   477 => x"85387184",
   478 => x"0752badc",
   479 => x"08802e85",
   480 => x"38719007",
   481 => x"5271bab0",
   482 => x"0c028805",
   483 => x"0d0402f4",
   484 => x"050d810b",
   485 => x"badc0c90",
   486 => x"5186932d",
   487 => x"810bfec4",
   488 => x"0c900bfe",
   489 => x"c00c840b",
   490 => x"fec40c83",
   491 => x"0bfecc0c",
   492 => x"a6f92da9",
   493 => x"8e2da6dc",
   494 => x"2da6dc2d",
   495 => x"81f82d81",
   496 => x"5184e62d",
   497 => x"a6dc2da6",
   498 => x"dc2d8151",
   499 => x"84e62db5",
   500 => x"c45185f2",
   501 => x"2d8452a0",
   502 => x"e72d92a6",
   503 => x"2dbab008",
   504 => x"802e8638",
   505 => x"fe528ff1",
   506 => x"04ff1252",
   507 => x"718024e7",
   508 => x"3871802e",
   509 => x"81833886",
   510 => x"c42db5dc",
   511 => x"5187b62d",
   512 => x"bab00880",
   513 => x"2e8f38b7",
   514 => x"a451ab91",
   515 => x"2d805184",
   516 => x"e62d909f",
   517 => x"04bab008",
   518 => x"518eb22d",
   519 => x"a99a2da7",
   520 => x"922dabaa",
   521 => x"2dbab008",
   522 => x"80c2d408",
   523 => x"882b80c2",
   524 => x"d80807fe",
   525 => x"d80c538e",
   526 => x"cf2dbab0",
   527 => x"08bad808",
   528 => x"2ea238ba",
   529 => x"b008bad8",
   530 => x"0cbab008",
   531 => x"fec00c84",
   532 => x"52725184",
   533 => x"e62da6dc",
   534 => x"2da6dc2d",
   535 => x"ff125271",
   536 => x"8025ee38",
   537 => x"72802e89",
   538 => x"388a0bfe",
   539 => x"c40c909f",
   540 => x"04820bfe",
   541 => x"c40c909f",
   542 => x"04b5e851",
   543 => x"85f22d80",
   544 => x"0bbab00c",
   545 => x"028c050d",
   546 => x"0402e805",
   547 => x"0d77797b",
   548 => x"58555580",
   549 => x"53727625",
   550 => x"a3387470",
   551 => x"81055680",
   552 => x"f52d7470",
   553 => x"81055680",
   554 => x"f52d5252",
   555 => x"71712e86",
   556 => x"38815191",
   557 => x"be048113",
   558 => x"53919504",
   559 => x"805170ba",
   560 => x"b00c0298",
   561 => x"050d0402",
   562 => x"f0050d75",
   563 => x"5372802e",
   564 => x"a2387280",
   565 => x"c2940c80",
   566 => x"c1e808fe",
   567 => x"14712980",
   568 => x"c1fc0805",
   569 => x"80c2980c",
   570 => x"70842b80",
   571 => x"c1f40c54",
   572 => x"92a10480",
   573 => x"c2800880",
   574 => x"c2940c80",
   575 => x"c2840880",
   576 => x"c2980c80",
   577 => x"c1f00880",
   578 => x"2e8b3880",
   579 => x"c1e80884",
   580 => x"2b53929c",
   581 => x"0480c288",
   582 => x"08842b53",
   583 => x"7280c1f4",
   584 => x"0c029005",
   585 => x"0d0402d8",
   586 => x"050d800b",
   587 => x"80c1f00c",
   588 => x"bde85280",
   589 => x"51a3d12d",
   590 => x"bab00854",
   591 => x"bab0088c",
   592 => x"38b5fc51",
   593 => x"85f22d73",
   594 => x"5597e804",
   595 => x"8056810b",
   596 => x"80c29c0c",
   597 => x"8853b688",
   598 => x"52be9e51",
   599 => x"91892dba",
   600 => x"b008762e",
   601 => x"09810688",
   602 => x"38bab008",
   603 => x"80c29c0c",
   604 => x"8853b694",
   605 => x"52beba51",
   606 => x"91892dba",
   607 => x"b0088838",
   608 => x"bab00880",
   609 => x"c29c0c80",
   610 => x"c29c0880",
   611 => x"2e80fc38",
   612 => x"80c1ae0b",
   613 => x"80f52d80",
   614 => x"c1af0b80",
   615 => x"f52d7198",
   616 => x"2b71902b",
   617 => x"0780c1b0",
   618 => x"0b80f52d",
   619 => x"70882b72",
   620 => x"0780c1b1",
   621 => x"0b80f52d",
   622 => x"710780c1",
   623 => x"e60b80f5",
   624 => x"2d80c1e7",
   625 => x"0b80f52d",
   626 => x"71882b07",
   627 => x"535f5452",
   628 => x"5a565755",
   629 => x"7381abaa",
   630 => x"2e098106",
   631 => x"8d387551",
   632 => x"a4f12dba",
   633 => x"b0085693",
   634 => x"f7047382",
   635 => x"d4d52e87",
   636 => x"38b6a051",
   637 => x"94b904bd",
   638 => x"e8527551",
   639 => x"a3d12dba",
   640 => x"b00855ba",
   641 => x"b008802e",
   642 => x"83de3888",
   643 => x"53b69452",
   644 => x"beba5191",
   645 => x"892dbab0",
   646 => x"088a3881",
   647 => x"0b80c1f0",
   648 => x"0c94bf04",
   649 => x"8853b688",
   650 => x"52be9e51",
   651 => x"91892dba",
   652 => x"b008802e",
   653 => x"8a38b6b4",
   654 => x"5185f22d",
   655 => x"959b0480",
   656 => x"c1e60b80",
   657 => x"f52d5473",
   658 => x"80d52e09",
   659 => x"810680cb",
   660 => x"3880c1e7",
   661 => x"0b80f52d",
   662 => x"547381aa",
   663 => x"2e098106",
   664 => x"ba38800b",
   665 => x"bde80b80",
   666 => x"f52d5654",
   667 => x"7481e92e",
   668 => x"83388154",
   669 => x"7481eb2e",
   670 => x"8c388055",
   671 => x"73752e09",
   672 => x"810682e4",
   673 => x"38bdf30b",
   674 => x"80f52d55",
   675 => x"748d38bd",
   676 => x"f40b80f5",
   677 => x"2d547382",
   678 => x"2e863880",
   679 => x"5597e804",
   680 => x"bdf50b80",
   681 => x"f52d7080",
   682 => x"c1e80cff",
   683 => x"0580c1ec",
   684 => x"0cbdf60b",
   685 => x"80f52dbd",
   686 => x"f70b80f5",
   687 => x"2d587605",
   688 => x"77828029",
   689 => x"057080c1",
   690 => x"f80cbdf8",
   691 => x"0b80f52d",
   692 => x"7080c28c",
   693 => x"0c80c1f0",
   694 => x"08595758",
   695 => x"76802e81",
   696 => x"ac388853",
   697 => x"b69452be",
   698 => x"ba519189",
   699 => x"2dbab008",
   700 => x"81f63880",
   701 => x"c1e80870",
   702 => x"842b80c1",
   703 => x"f40c7080",
   704 => x"c2880cbe",
   705 => x"8d0b80f5",
   706 => x"2dbe8c0b",
   707 => x"80f52d71",
   708 => x"82802905",
   709 => x"be8e0b80",
   710 => x"f52d7084",
   711 => x"80802912",
   712 => x"be8f0b80",
   713 => x"f52d7081",
   714 => x"800a2912",
   715 => x"7080c290",
   716 => x"0c80c28c",
   717 => x"08712980",
   718 => x"c1f80805",
   719 => x"7080c1fc",
   720 => x"0cbe950b",
   721 => x"80f52dbe",
   722 => x"940b80f5",
   723 => x"2d718280",
   724 => x"2905be96",
   725 => x"0b80f52d",
   726 => x"70848080",
   727 => x"2912be97",
   728 => x"0b80f52d",
   729 => x"70982b81",
   730 => x"f00a0672",
   731 => x"057080c2",
   732 => x"800cfe11",
   733 => x"7e297705",
   734 => x"80c2840c",
   735 => x"52595243",
   736 => x"545e5152",
   737 => x"59525d57",
   738 => x"595797e1",
   739 => x"04bdfa0b",
   740 => x"80f52dbd",
   741 => x"f90b80f5",
   742 => x"2d718280",
   743 => x"29057080",
   744 => x"c1f40c70",
   745 => x"a02983ff",
   746 => x"0570892a",
   747 => x"7080c288",
   748 => x"0cbdff0b",
   749 => x"80f52dbd",
   750 => x"fe0b80f5",
   751 => x"2d718280",
   752 => x"29057080",
   753 => x"c2900c7b",
   754 => x"71291e70",
   755 => x"80c2840c",
   756 => x"7d80c280",
   757 => x"0c730580",
   758 => x"c1fc0c55",
   759 => x"5e515155",
   760 => x"55805191",
   761 => x"c72d8155",
   762 => x"74bab00c",
   763 => x"02a8050d",
   764 => x"0402ec05",
   765 => x"0d767087",
   766 => x"2c7180ff",
   767 => x"06555654",
   768 => x"80c1f008",
   769 => x"8a387388",
   770 => x"2c7481ff",
   771 => x"065455bd",
   772 => x"e85280c1",
   773 => x"f8081551",
   774 => x"a3d12dba",
   775 => x"b00854ba",
   776 => x"b008802e",
   777 => x"b43880c1",
   778 => x"f008802e",
   779 => x"98387284",
   780 => x"29bde805",
   781 => x"70085253",
   782 => x"a4f12dba",
   783 => x"b008f00a",
   784 => x"065398d7",
   785 => x"047210bd",
   786 => x"e8057080",
   787 => x"e02d5253",
   788 => x"a5a12dba",
   789 => x"b0085372",
   790 => x"5473bab0",
   791 => x"0c029405",
   792 => x"0d0402ec",
   793 => x"050d7670",
   794 => x"842c80c2",
   795 => x"98080571",
   796 => x"8f065255",
   797 => x"53728938",
   798 => x"bde85273",
   799 => x"51a3d12d",
   800 => x"72a029bd",
   801 => x"e8055580",
   802 => x"7580f52d",
   803 => x"55537373",
   804 => x"2e833881",
   805 => x"537381e5",
   806 => x"2e9b3872",
   807 => x"802e9638",
   808 => x"8b1580f5",
   809 => x"2d70832a",
   810 => x"70810677",
   811 => x"53515454",
   812 => x"72802e83",
   813 => x"38805473",
   814 => x"bab00c02",
   815 => x"94050d04",
   816 => x"02cc050d",
   817 => x"7e605e5a",
   818 => x"800b80c2",
   819 => x"940880c2",
   820 => x"9808595c",
   821 => x"56805880",
   822 => x"c1f40878",
   823 => x"2e81b038",
   824 => x"778f06a0",
   825 => x"17575473",
   826 => x"8f38bde8",
   827 => x"52765181",
   828 => x"1757a3d1",
   829 => x"2dbde856",
   830 => x"807680f5",
   831 => x"2d565474",
   832 => x"742e8338",
   833 => x"81547481",
   834 => x"e52e80f7",
   835 => x"38817075",
   836 => x"06555c73",
   837 => x"802e80eb",
   838 => x"388b1680",
   839 => x"f52d9806",
   840 => x"597880df",
   841 => x"388b537c",
   842 => x"52755191",
   843 => x"892dbab0",
   844 => x"0880d038",
   845 => x"9c160851",
   846 => x"a4f12dba",
   847 => x"b008841b",
   848 => x"0c9a1680",
   849 => x"e02d51a5",
   850 => x"a12dbab0",
   851 => x"08bab008",
   852 => x"881c0cba",
   853 => x"b0085555",
   854 => x"80c1f008",
   855 => x"802e9838",
   856 => x"941680e0",
   857 => x"2d51a5a1",
   858 => x"2dbab008",
   859 => x"902b83ff",
   860 => x"f00a0670",
   861 => x"16515473",
   862 => x"881b0c78",
   863 => x"7a0c7b54",
   864 => x"9bc80481",
   865 => x"185880c1",
   866 => x"f4087826",
   867 => x"fed23880",
   868 => x"c1f00880",
   869 => x"2eb0387a",
   870 => x"5197f12d",
   871 => x"bab008ba",
   872 => x"b00880ff",
   873 => x"fffff806",
   874 => x"555b7380",
   875 => x"fffffff8",
   876 => x"2e9438ba",
   877 => x"b008fe05",
   878 => x"80c1e808",
   879 => x"2980c1fc",
   880 => x"08055799",
   881 => x"d5048054",
   882 => x"73bab00c",
   883 => x"02b4050d",
   884 => x"0402f405",
   885 => x"0d747008",
   886 => x"8105710c",
   887 => x"700880c1",
   888 => x"ec080653",
   889 => x"53718e38",
   890 => x"88130851",
   891 => x"97f12dba",
   892 => x"b0088814",
   893 => x"0c810bba",
   894 => x"b00c028c",
   895 => x"050d0402",
   896 => x"f0050d75",
   897 => x"881108fe",
   898 => x"0580c1e8",
   899 => x"082980c1",
   900 => x"fc081172",
   901 => x"0880c1ec",
   902 => x"08060579",
   903 => x"55535454",
   904 => x"a3d12d02",
   905 => x"90050d04",
   906 => x"02f0050d",
   907 => x"75881108",
   908 => x"fe0580c1",
   909 => x"e8082980",
   910 => x"c1fc0811",
   911 => x"720880c1",
   912 => x"ec080605",
   913 => x"79555354",
   914 => x"54a2912d",
   915 => x"0290050d",
   916 => x"0480c1f0",
   917 => x"08bab00c",
   918 => x"0402f405",
   919 => x"0dd45281",
   920 => x"ff720c71",
   921 => x"085381ff",
   922 => x"720c7288",
   923 => x"2b83fe80",
   924 => x"06720870",
   925 => x"81ff0651",
   926 => x"525381ff",
   927 => x"720c7271",
   928 => x"07882b72",
   929 => x"087081ff",
   930 => x"06515253",
   931 => x"81ff720c",
   932 => x"72710788",
   933 => x"2b720870",
   934 => x"81ff0672",
   935 => x"07bab00c",
   936 => x"5253028c",
   937 => x"050d0402",
   938 => x"f4050d74",
   939 => x"767181ff",
   940 => x"06d40c53",
   941 => x"5380c2a0",
   942 => x"08853871",
   943 => x"892b5271",
   944 => x"982ad40c",
   945 => x"71902a70",
   946 => x"81ff06d4",
   947 => x"0c517188",
   948 => x"2a7081ff",
   949 => x"06d40c51",
   950 => x"7181ff06",
   951 => x"d40c7290",
   952 => x"2a7081ff",
   953 => x"06d40c51",
   954 => x"d4087081",
   955 => x"ff065151",
   956 => x"82b8bf52",
   957 => x"7081ff2e",
   958 => x"09810694",
   959 => x"3881ff0b",
   960 => x"d40cd408",
   961 => x"7081ff06",
   962 => x"ff145451",
   963 => x"5171e538",
   964 => x"70bab00c",
   965 => x"028c050d",
   966 => x"0402fc05",
   967 => x"0d81c751",
   968 => x"81ff0bd4",
   969 => x"0cff1151",
   970 => x"708025f4",
   971 => x"38028405",
   972 => x"0d0402f0",
   973 => x"050d9e99",
   974 => x"2d8fcf53",
   975 => x"805287fc",
   976 => x"80f7519d",
   977 => x"a72dbab0",
   978 => x"0854bab0",
   979 => x"08812e09",
   980 => x"8106a338",
   981 => x"81ff0bd4",
   982 => x"0c820a52",
   983 => x"849c80e9",
   984 => x"519da72d",
   985 => x"bab0088b",
   986 => x"3881ff0b",
   987 => x"d40c7353",
   988 => x"9efc049e",
   989 => x"992dff13",
   990 => x"5372c138",
   991 => x"72bab00c",
   992 => x"0290050d",
   993 => x"0402f405",
   994 => x"0d81ff0b",
   995 => x"d40c9353",
   996 => x"805287fc",
   997 => x"80c1519d",
   998 => x"a72dbab0",
   999 => x"088b3881",
  1000 => x"ff0bd40c",
  1001 => x"81539fb2",
  1002 => x"049e992d",
  1003 => x"ff135372",
  1004 => x"df3872ba",
  1005 => x"b00c028c",
  1006 => x"050d0402",
  1007 => x"f0050d9e",
  1008 => x"992d83aa",
  1009 => x"52849c80",
  1010 => x"c8519da7",
  1011 => x"2dbab008",
  1012 => x"812e0981",
  1013 => x"0692389c",
  1014 => x"d92dbab0",
  1015 => x"0883ffff",
  1016 => x"06537283",
  1017 => x"aa2e9738",
  1018 => x"9f852d9f",
  1019 => x"f9048154",
  1020 => x"a0de04b6",
  1021 => x"c05185f2",
  1022 => x"2d8054a0",
  1023 => x"de0481ff",
  1024 => x"0bd40cb1",
  1025 => x"539eb22d",
  1026 => x"bab00880",
  1027 => x"2e80c038",
  1028 => x"805287fc",
  1029 => x"80fa519d",
  1030 => x"a72dbab0",
  1031 => x"08b13881",
  1032 => x"ff0bd40c",
  1033 => x"d4085381",
  1034 => x"ff0bd40c",
  1035 => x"81ff0bd4",
  1036 => x"0c81ff0b",
  1037 => x"d40c81ff",
  1038 => x"0bd40c72",
  1039 => x"862a7081",
  1040 => x"06bab008",
  1041 => x"56515372",
  1042 => x"802e9338",
  1043 => x"9fee0472",
  1044 => x"822eff9f",
  1045 => x"38ff1353",
  1046 => x"72ffaa38",
  1047 => x"725473ba",
  1048 => x"b00c0290",
  1049 => x"050d0402",
  1050 => x"f0050d81",
  1051 => x"0b80c2a0",
  1052 => x"0c8454d0",
  1053 => x"08708f2a",
  1054 => x"70810651",
  1055 => x"515372f3",
  1056 => x"3872d00c",
  1057 => x"9e992db6",
  1058 => x"d05185f2",
  1059 => x"2dd00870",
  1060 => x"8f2a7081",
  1061 => x"06515153",
  1062 => x"72f33881",
  1063 => x"0bd00cb1",
  1064 => x"53805284",
  1065 => x"d480c051",
  1066 => x"9da72dba",
  1067 => x"b008812e",
  1068 => x"a1387282",
  1069 => x"2e098106",
  1070 => x"8c38b6dc",
  1071 => x"5185f22d",
  1072 => x"8053a288",
  1073 => x"04ff1353",
  1074 => x"72d738ff",
  1075 => x"145473ff",
  1076 => x"a2389fbb",
  1077 => x"2dbab008",
  1078 => x"80c2a00c",
  1079 => x"bab0088b",
  1080 => x"38815287",
  1081 => x"fc80d051",
  1082 => x"9da72d81",
  1083 => x"ff0bd40c",
  1084 => x"d008708f",
  1085 => x"2a708106",
  1086 => x"51515372",
  1087 => x"f33872d0",
  1088 => x"0c81ff0b",
  1089 => x"d40c8153",
  1090 => x"72bab00c",
  1091 => x"0290050d",
  1092 => x"0402e805",
  1093 => x"0d785681",
  1094 => x"ff0bd40c",
  1095 => x"d008708f",
  1096 => x"2a708106",
  1097 => x"51515372",
  1098 => x"f3388281",
  1099 => x"0bd00c81",
  1100 => x"ff0bd40c",
  1101 => x"775287fc",
  1102 => x"80d8519d",
  1103 => x"a72dbab0",
  1104 => x"08802e8c",
  1105 => x"38b6f451",
  1106 => x"85f22d81",
  1107 => x"53a3c804",
  1108 => x"81ff0bd4",
  1109 => x"0c81fe0b",
  1110 => x"d40c80ff",
  1111 => x"55757084",
  1112 => x"05570870",
  1113 => x"982ad40c",
  1114 => x"70902c70",
  1115 => x"81ff06d4",
  1116 => x"0c547088",
  1117 => x"2c7081ff",
  1118 => x"06d40c54",
  1119 => x"7081ff06",
  1120 => x"d40c54ff",
  1121 => x"15557480",
  1122 => x"25d33881",
  1123 => x"ff0bd40c",
  1124 => x"81ff0bd4",
  1125 => x"0c81ff0b",
  1126 => x"d40c868d",
  1127 => x"a05481ff",
  1128 => x"0bd40cd4",
  1129 => x"0881ff06",
  1130 => x"55748738",
  1131 => x"ff145473",
  1132 => x"ed3881ff",
  1133 => x"0bd40cd0",
  1134 => x"08708f2a",
  1135 => x"70810651",
  1136 => x"515372f3",
  1137 => x"3872d00c",
  1138 => x"72bab00c",
  1139 => x"0298050d",
  1140 => x"0402e805",
  1141 => x"0d785580",
  1142 => x"5681ff0b",
  1143 => x"d40cd008",
  1144 => x"708f2a70",
  1145 => x"81065151",
  1146 => x"5372f338",
  1147 => x"82810bd0",
  1148 => x"0c81ff0b",
  1149 => x"d40c7752",
  1150 => x"87fc80d1",
  1151 => x"519da72d",
  1152 => x"80dbc6df",
  1153 => x"54bab008",
  1154 => x"802e8a38",
  1155 => x"b7845185",
  1156 => x"f22da4e8",
  1157 => x"0481ff0b",
  1158 => x"d40cd408",
  1159 => x"7081ff06",
  1160 => x"51537281",
  1161 => x"fe2e0981",
  1162 => x"069d3880",
  1163 => x"ff539cd9",
  1164 => x"2dbab008",
  1165 => x"75708405",
  1166 => x"570cff13",
  1167 => x"53728025",
  1168 => x"ed388156",
  1169 => x"a4cd04ff",
  1170 => x"145473c9",
  1171 => x"3881ff0b",
  1172 => x"d40c81ff",
  1173 => x"0bd40cd0",
  1174 => x"08708f2a",
  1175 => x"70810651",
  1176 => x"515372f3",
  1177 => x"3872d00c",
  1178 => x"75bab00c",
  1179 => x"0298050d",
  1180 => x"0402f405",
  1181 => x"0d747088",
  1182 => x"2a83fe80",
  1183 => x"06707298",
  1184 => x"2a077288",
  1185 => x"2b87fc80",
  1186 => x"80067398",
  1187 => x"2b81f00a",
  1188 => x"06717307",
  1189 => x"07bab00c",
  1190 => x"56515351",
  1191 => x"028c050d",
  1192 => x"0402f805",
  1193 => x"0d028e05",
  1194 => x"80f52d74",
  1195 => x"882b0770",
  1196 => x"83ffff06",
  1197 => x"bab00c51",
  1198 => x"0288050d",
  1199 => x"0402fc05",
  1200 => x"0d725180",
  1201 => x"710c800b",
  1202 => x"84120c02",
  1203 => x"84050d04",
  1204 => x"02f0050d",
  1205 => x"75700884",
  1206 => x"12085353",
  1207 => x"53ff5471",
  1208 => x"712ea838",
  1209 => x"a9942d84",
  1210 => x"13087084",
  1211 => x"29148811",
  1212 => x"70087081",
  1213 => x"ff068418",
  1214 => x"08811187",
  1215 => x"06841a0c",
  1216 => x"53515551",
  1217 => x"5151a98e",
  1218 => x"2d715473",
  1219 => x"bab00c02",
  1220 => x"90050d04",
  1221 => x"02f8050d",
  1222 => x"a9942de0",
  1223 => x"08708b2a",
  1224 => x"70810651",
  1225 => x"52527080",
  1226 => x"2ea13880",
  1227 => x"c2a40870",
  1228 => x"842980c2",
  1229 => x"ac057381",
  1230 => x"ff06710c",
  1231 => x"515180c2",
  1232 => x"a4088111",
  1233 => x"870680c2",
  1234 => x"a40c5180",
  1235 => x"0b80c2cc",
  1236 => x"0ca9872d",
  1237 => x"a98e2d02",
  1238 => x"88050d04",
  1239 => x"02fc050d",
  1240 => x"a9942d81",
  1241 => x"0b80c2cc",
  1242 => x"0ca98e2d",
  1243 => x"80c2cc08",
  1244 => x"5170f938",
  1245 => x"0284050d",
  1246 => x"0402fc05",
  1247 => x"0d80c2a4",
  1248 => x"51a5bd2d",
  1249 => x"a69451a9",
  1250 => x"832da8ad",
  1251 => x"2d028405",
  1252 => x"0d0402f4",
  1253 => x"050da894",
  1254 => x"04bab008",
  1255 => x"81f02e09",
  1256 => x"81068938",
  1257 => x"810bbaa4",
  1258 => x"0ca89404",
  1259 => x"bab00881",
  1260 => x"e02e0981",
  1261 => x"06893881",
  1262 => x"0bbaa80c",
  1263 => x"a89404ba",
  1264 => x"b00852ba",
  1265 => x"a808802e",
  1266 => x"8838bab0",
  1267 => x"08818005",
  1268 => x"5271842c",
  1269 => x"728f0653",
  1270 => x"53baa408",
  1271 => x"802e9938",
  1272 => x"728429b9",
  1273 => x"e4057213",
  1274 => x"81712b70",
  1275 => x"09730806",
  1276 => x"730c5153",
  1277 => x"53a88a04",
  1278 => x"728429b9",
  1279 => x"e4057213",
  1280 => x"83712b72",
  1281 => x"0807720c",
  1282 => x"5353800b",
  1283 => x"baa80c80",
  1284 => x"0bbaa40c",
  1285 => x"80c2a451",
  1286 => x"a5d02dba",
  1287 => x"b008ff24",
  1288 => x"fef73880",
  1289 => x"0bbab00c",
  1290 => x"028c050d",
  1291 => x"0402f805",
  1292 => x"0db9e452",
  1293 => x"8f518072",
  1294 => x"70840554",
  1295 => x"0cff1151",
  1296 => x"708025f2",
  1297 => x"38028805",
  1298 => x"0d0402f0",
  1299 => x"050d7551",
  1300 => x"a9942d70",
  1301 => x"822cfc06",
  1302 => x"b9e41172",
  1303 => x"109e0671",
  1304 => x"0870722a",
  1305 => x"70830682",
  1306 => x"742b7009",
  1307 => x"7406760c",
  1308 => x"54515657",
  1309 => x"535153a9",
  1310 => x"8e2d71ba",
  1311 => x"b00c0290",
  1312 => x"050d0471",
  1313 => x"980c04ff",
  1314 => x"b008bab0",
  1315 => x"0c04810b",
  1316 => x"ffb00c04",
  1317 => x"800bffb0",
  1318 => x"0c0402fc",
  1319 => x"050d810b",
  1320 => x"baac0c81",
  1321 => x"5184e62d",
  1322 => x"0284050d",
  1323 => x"0402fc05",
  1324 => x"0d800bba",
  1325 => x"ac0c8051",
  1326 => x"84e62d02",
  1327 => x"84050d04",
  1328 => x"02ec050d",
  1329 => x"76548052",
  1330 => x"870b8815",
  1331 => x"80f52d56",
  1332 => x"53747224",
  1333 => x"8338a053",
  1334 => x"725182ef",
  1335 => x"2d81128b",
  1336 => x"1580f52d",
  1337 => x"54527272",
  1338 => x"25de3802",
  1339 => x"94050d04",
  1340 => x"02f0050d",
  1341 => x"80c2dc08",
  1342 => x"5481f82d",
  1343 => x"800b80c2",
  1344 => x"e00c7308",
  1345 => x"802e8184",
  1346 => x"38820bba",
  1347 => x"c40c80c2",
  1348 => x"e0088f06",
  1349 => x"bac00c73",
  1350 => x"08527183",
  1351 => x"2e963871",
  1352 => x"83268938",
  1353 => x"71812eaf",
  1354 => x"38aaf504",
  1355 => x"71852e9f",
  1356 => x"38aaf504",
  1357 => x"881480f5",
  1358 => x"2d841508",
  1359 => x"b7945354",
  1360 => x"5285f22d",
  1361 => x"71842913",
  1362 => x"70085252",
  1363 => x"aaf90473",
  1364 => x"51a9c02d",
  1365 => x"aaf50480",
  1366 => x"c2d00888",
  1367 => x"15082c70",
  1368 => x"81065152",
  1369 => x"71802e87",
  1370 => x"38b79851",
  1371 => x"aaf204b7",
  1372 => x"9c5185f2",
  1373 => x"2d841408",
  1374 => x"5185f22d",
  1375 => x"80c2e008",
  1376 => x"810580c2",
  1377 => x"e00c8c14",
  1378 => x"54aa8204",
  1379 => x"0290050d",
  1380 => x"047180c2",
  1381 => x"dc0ca9f0",
  1382 => x"2d80c2e0",
  1383 => x"08ff0580",
  1384 => x"c2e40c04",
  1385 => x"7180c2e8",
  1386 => x"0c0402e8",
  1387 => x"050d80c2",
  1388 => x"dc0880c2",
  1389 => x"e8085755",
  1390 => x"80f851a8",
  1391 => x"ca2dbab0",
  1392 => x"08812a70",
  1393 => x"81065152",
  1394 => x"719b3887",
  1395 => x"51a8ca2d",
  1396 => x"bab00881",
  1397 => x"2a708106",
  1398 => x"51527180",
  1399 => x"2eb138ab",
  1400 => x"e504a792",
  1401 => x"2d8751a8",
  1402 => x"ca2dbab0",
  1403 => x"08f438ab",
  1404 => x"f504a792",
  1405 => x"2d80f851",
  1406 => x"a8ca2dba",
  1407 => x"b008f338",
  1408 => x"baac0881",
  1409 => x"3270baac",
  1410 => x"0c705252",
  1411 => x"84e62d80",
  1412 => x"0b80c2d4",
  1413 => x"0c800b80",
  1414 => x"c2d80cba",
  1415 => x"ac0882fd",
  1416 => x"3880da51",
  1417 => x"a8ca2dba",
  1418 => x"b008802e",
  1419 => x"8c3880c2",
  1420 => x"d4088180",
  1421 => x"0780c2d4",
  1422 => x"0c80d951",
  1423 => x"a8ca2dba",
  1424 => x"b008802e",
  1425 => x"8c3880c2",
  1426 => x"d40880c0",
  1427 => x"0780c2d4",
  1428 => x"0c819451",
  1429 => x"a8ca2dba",
  1430 => x"b008802e",
  1431 => x"8b3880c2",
  1432 => x"d4089007",
  1433 => x"80c2d40c",
  1434 => x"819151a8",
  1435 => x"ca2dbab0",
  1436 => x"08802e8b",
  1437 => x"3880c2d4",
  1438 => x"08a00780",
  1439 => x"c2d40c81",
  1440 => x"f551a8ca",
  1441 => x"2dbab008",
  1442 => x"802e8b38",
  1443 => x"80c2d408",
  1444 => x"810780c2",
  1445 => x"d40c81f2",
  1446 => x"51a8ca2d",
  1447 => x"bab00880",
  1448 => x"2e8b3880",
  1449 => x"c2d40882",
  1450 => x"0780c2d4",
  1451 => x"0c81eb51",
  1452 => x"a8ca2dba",
  1453 => x"b008802e",
  1454 => x"8b3880c2",
  1455 => x"d4088407",
  1456 => x"80c2d40c",
  1457 => x"81f451a8",
  1458 => x"ca2dbab0",
  1459 => x"08802e8b",
  1460 => x"3880c2d4",
  1461 => x"08880780",
  1462 => x"c2d40c80",
  1463 => x"d851a8ca",
  1464 => x"2dbab008",
  1465 => x"802e8c38",
  1466 => x"80c2d808",
  1467 => x"81800780",
  1468 => x"c2d80c92",
  1469 => x"51a8ca2d",
  1470 => x"bab00880",
  1471 => x"2e8c3880",
  1472 => x"c2d80880",
  1473 => x"c00780c2",
  1474 => x"d80c9451",
  1475 => x"a8ca2dba",
  1476 => x"b008802e",
  1477 => x"8b3880c2",
  1478 => x"d8089007",
  1479 => x"80c2d80c",
  1480 => x"9151a8ca",
  1481 => x"2dbab008",
  1482 => x"802e8b38",
  1483 => x"80c2d808",
  1484 => x"a00780c2",
  1485 => x"d80c9d51",
  1486 => x"a8ca2dba",
  1487 => x"b008802e",
  1488 => x"8b3880c2",
  1489 => x"d8088107",
  1490 => x"80c2d80c",
  1491 => x"9b51a8ca",
  1492 => x"2dbab008",
  1493 => x"802e8b38",
  1494 => x"80c2d808",
  1495 => x"820780c2",
  1496 => x"d80c9c51",
  1497 => x"a8ca2dba",
  1498 => x"b008802e",
  1499 => x"8b3880c2",
  1500 => x"d8088407",
  1501 => x"80c2d80c",
  1502 => x"a351a8ca",
  1503 => x"2dbab008",
  1504 => x"802e8b38",
  1505 => x"80c2d808",
  1506 => x"880780c2",
  1507 => x"d80c81fd",
  1508 => x"51a8ca2d",
  1509 => x"81fa51a8",
  1510 => x"ca2db495",
  1511 => x"0481f551",
  1512 => x"a8ca2dba",
  1513 => x"b008812a",
  1514 => x"70810651",
  1515 => x"5271802e",
  1516 => x"b33880c2",
  1517 => x"e4085271",
  1518 => x"802e8a38",
  1519 => x"ff1280c2",
  1520 => x"e40cafe4",
  1521 => x"0480c2e0",
  1522 => x"081080c2",
  1523 => x"e0080570",
  1524 => x"84291651",
  1525 => x"52881208",
  1526 => x"802e8938",
  1527 => x"ff518812",
  1528 => x"0852712d",
  1529 => x"81f251a8",
  1530 => x"ca2dbab0",
  1531 => x"08812a70",
  1532 => x"81065152",
  1533 => x"71802eb4",
  1534 => x"3880c2e0",
  1535 => x"08ff1180",
  1536 => x"c2e40856",
  1537 => x"53537372",
  1538 => x"258a3881",
  1539 => x"1480c2e4",
  1540 => x"0cb0ac04",
  1541 => x"72101370",
  1542 => x"84291651",
  1543 => x"52881208",
  1544 => x"802e8938",
  1545 => x"fe518812",
  1546 => x"0852712d",
  1547 => x"81fd51a8",
  1548 => x"ca2dbab0",
  1549 => x"08812a70",
  1550 => x"81065152",
  1551 => x"71802e87",
  1552 => x"38800b80",
  1553 => x"c2e40c81",
  1554 => x"fa51a8ca",
  1555 => x"2dbab008",
  1556 => x"812a7081",
  1557 => x"06515271",
  1558 => x"802e8b38",
  1559 => x"80c2e008",
  1560 => x"ff0580c2",
  1561 => x"e40c80c2",
  1562 => x"e4087053",
  1563 => x"5473802e",
  1564 => x"8a388c15",
  1565 => x"ff155555",
  1566 => x"b0ed0482",
  1567 => x"0bbac40c",
  1568 => x"718f06ba",
  1569 => x"c00c81eb",
  1570 => x"51a8ca2d",
  1571 => x"bab00881",
  1572 => x"2a708106",
  1573 => x"51527180",
  1574 => x"2ead3874",
  1575 => x"08852e09",
  1576 => x"8106a438",
  1577 => x"881580f5",
  1578 => x"2dff0552",
  1579 => x"71881681",
  1580 => x"b72d7198",
  1581 => x"2b527180",
  1582 => x"25883880",
  1583 => x"0b881681",
  1584 => x"b72d7451",
  1585 => x"a9c02d81",
  1586 => x"f451a8ca",
  1587 => x"2dbab008",
  1588 => x"812a7081",
  1589 => x"06515271",
  1590 => x"802eb338",
  1591 => x"7408852e",
  1592 => x"098106aa",
  1593 => x"38881580",
  1594 => x"f52d8105",
  1595 => x"52718816",
  1596 => x"81b72d71",
  1597 => x"81ff068b",
  1598 => x"1680f52d",
  1599 => x"54527272",
  1600 => x"27873872",
  1601 => x"881681b7",
  1602 => x"2d7451a9",
  1603 => x"c02d80da",
  1604 => x"51a8ca2d",
  1605 => x"bab00881",
  1606 => x"2a708106",
  1607 => x"51527180",
  1608 => x"2e81ac38",
  1609 => x"80c2dc08",
  1610 => x"80c2e408",
  1611 => x"55537380",
  1612 => x"2e8a388c",
  1613 => x"13ff1555",
  1614 => x"53b2ae04",
  1615 => x"72085271",
  1616 => x"822ea638",
  1617 => x"71822689",
  1618 => x"3871812e",
  1619 => x"aa38b3cf",
  1620 => x"0471832e",
  1621 => x"b4387184",
  1622 => x"2e098106",
  1623 => x"80f13888",
  1624 => x"130851ab",
  1625 => x"912db3cf",
  1626 => x"0480c2e4",
  1627 => x"08518813",
  1628 => x"0852712d",
  1629 => x"b3cf0481",
  1630 => x"0b881408",
  1631 => x"2b80c2d0",
  1632 => x"083280c2",
  1633 => x"d00cb3a4",
  1634 => x"04881380",
  1635 => x"f52d8105",
  1636 => x"8b1480f5",
  1637 => x"2d535471",
  1638 => x"74248338",
  1639 => x"80547388",
  1640 => x"1481b72d",
  1641 => x"a9f02db3",
  1642 => x"cf047508",
  1643 => x"802ea338",
  1644 => x"750851a8",
  1645 => x"ca2dbab0",
  1646 => x"08810652",
  1647 => x"71802e8c",
  1648 => x"3880c2e4",
  1649 => x"08518416",
  1650 => x"0852712d",
  1651 => x"88165675",
  1652 => x"d9388054",
  1653 => x"800bbac4",
  1654 => x"0c738f06",
  1655 => x"bac00ca0",
  1656 => x"527380c2",
  1657 => x"e4082e09",
  1658 => x"81069938",
  1659 => x"80c2e008",
  1660 => x"ff057432",
  1661 => x"70098105",
  1662 => x"7072079f",
  1663 => x"2a917131",
  1664 => x"51515353",
  1665 => x"715182ef",
  1666 => x"2d811454",
  1667 => x"8e7425c4",
  1668 => x"38baac08",
  1669 => x"5271bab0",
  1670 => x"0c029805",
  1671 => x"0d040000",
  1672 => x"00ffffff",
  1673 => x"ff00ffff",
  1674 => x"ffff00ff",
  1675 => x"ffffff00",
  1676 => x"52657365",
  1677 => x"74000000",
  1678 => x"53617665",
  1679 => x"20736574",
  1680 => x"74696e67",
  1681 => x"73000000",
  1682 => x"5363616e",
  1683 => x"6c696e65",
  1684 => x"73000000",
  1685 => x"4c6f6164",
  1686 => x"20524f4d",
  1687 => x"20100000",
  1688 => x"45786974",
  1689 => x"00000000",
  1690 => x"50432045",
  1691 => x"6e67696e",
  1692 => x"65206d6f",
  1693 => x"64650000",
  1694 => x"54757262",
  1695 => x"6f677261",
  1696 => x"66782031",
  1697 => x"36206d6f",
  1698 => x"64650000",
  1699 => x"56474120",
  1700 => x"2d203331",
  1701 => x"4b487a2c",
  1702 => x"20363048",
  1703 => x"7a000000",
  1704 => x"5456202d",
  1705 => x"20343830",
  1706 => x"692c2036",
  1707 => x"30487a00",
  1708 => x"4261636b",
  1709 => x"00000000",
  1710 => x"46504741",
  1711 => x"50434520",
  1712 => x"43464700",
  1713 => x"496e6974",
  1714 => x"69616c69",
  1715 => x"7a696e67",
  1716 => x"20534420",
  1717 => x"63617264",
  1718 => x"0a000000",
  1719 => x"424f4f54",
  1720 => x"20202020",
  1721 => x"50434500",
  1722 => x"43617264",
  1723 => x"20696e69",
  1724 => x"74206661",
  1725 => x"696c6564",
  1726 => x"0a000000",
  1727 => x"4d425220",
  1728 => x"6661696c",
  1729 => x"0a000000",
  1730 => x"46415431",
  1731 => x"36202020",
  1732 => x"00000000",
  1733 => x"46415433",
  1734 => x"32202020",
  1735 => x"00000000",
  1736 => x"4e6f2070",
  1737 => x"61727469",
  1738 => x"74696f6e",
  1739 => x"20736967",
  1740 => x"0a000000",
  1741 => x"42616420",
  1742 => x"70617274",
  1743 => x"0a000000",
  1744 => x"53444843",
  1745 => x"20657272",
  1746 => x"6f72210a",
  1747 => x"00000000",
  1748 => x"53442069",
  1749 => x"6e69742e",
  1750 => x"2e2e0a00",
  1751 => x"53442063",
  1752 => x"61726420",
  1753 => x"72657365",
  1754 => x"74206661",
  1755 => x"696c6564",
  1756 => x"210a0000",
  1757 => x"57726974",
  1758 => x"65206661",
  1759 => x"696c6564",
  1760 => x"0a000000",
  1761 => x"52656164",
  1762 => x"20666169",
  1763 => x"6c65640a",
  1764 => x"00000000",
  1765 => x"16200000",
  1766 => x"14200000",
  1767 => x"15200000",
  1768 => x"00000002",
  1769 => x"00000002",
  1770 => x"00001a30",
  1771 => x"000004b2",
  1772 => x"00000002",
  1773 => x"00001a38",
  1774 => x"00000379",
  1775 => x"00000003",
  1776 => x"00001c0c",
  1777 => x"00000002",
  1778 => x"00000001",
  1779 => x"00001a48",
  1780 => x"00000001",
  1781 => x"00000003",
  1782 => x"00001c04",
  1783 => x"00000002",
  1784 => x"00000002",
  1785 => x"00001a54",
  1786 => x"00000732",
  1787 => x"00000002",
  1788 => x"00001a60",
  1789 => x"000014ad",
  1790 => x"00000000",
  1791 => x"00000000",
  1792 => x"00000000",
  1793 => x"00001a68",
  1794 => x"00001a78",
  1795 => x"00001a8c",
  1796 => x"00001aa0",
  1797 => x"0000004d",
  1798 => x"00000706",
  1799 => x"0000002c",
  1800 => x"0000071c",
  1801 => x"00000000",
  1802 => x"00000000",
  1803 => x"00000002",
  1804 => x"00001d60",
  1805 => x"000004c7",
  1806 => x"00000002",
  1807 => x"00001d7e",
  1808 => x"000004c7",
  1809 => x"00000002",
  1810 => x"00001d9c",
  1811 => x"000004c7",
  1812 => x"00000002",
  1813 => x"00001dba",
  1814 => x"000004c7",
  1815 => x"00000002",
  1816 => x"00001dd8",
  1817 => x"000004c7",
  1818 => x"00000002",
  1819 => x"00001df6",
  1820 => x"000004c7",
  1821 => x"00000002",
  1822 => x"00001e14",
  1823 => x"000004c7",
  1824 => x"00000002",
  1825 => x"00001e32",
  1826 => x"000004c7",
  1827 => x"00000002",
  1828 => x"00001e50",
  1829 => x"000004c7",
  1830 => x"00000002",
  1831 => x"00001e6e",
  1832 => x"000004c7",
  1833 => x"00000002",
  1834 => x"00001e8c",
  1835 => x"000004c7",
  1836 => x"00000002",
  1837 => x"00001eaa",
  1838 => x"000004c7",
  1839 => x"00000002",
  1840 => x"00001ec8",
  1841 => x"000004c7",
  1842 => x"00000004",
  1843 => x"00001ab0",
  1844 => x"00001ba4",
  1845 => x"00000000",
  1846 => x"00000000",
  1847 => x"0000069a",
  1848 => x"00000000",
  1849 => x"00000000",
  1850 => x"00000000",
  1851 => x"00000000",
  1852 => x"00000000",
  1853 => x"00000000",
  1854 => x"00000000",
  1855 => x"00000000",
  1856 => x"00000000",
  1857 => x"00000000",
  1858 => x"00000000",
  1859 => x"00000000",
  1860 => x"00000000",
  1861 => x"00000000",
  1862 => x"00000000",
  1863 => x"00000000",
  1864 => x"00000000",
  1865 => x"00000000",
  1866 => x"00000000",
  1867 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

