-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bac",
     9 => x"f0080b0b",
    10 => x"0bacf408",
    11 => x"0b0b0bac",
    12 => x"f8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"acf80c0b",
    16 => x"0b0bacf4",
    17 => x"0c0b0b0b",
    18 => x"acf00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba8bc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"acf070b2",
    57 => x"8c278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8ab10402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"ad800c9f",
    65 => x"0bad840c",
    66 => x"a0717081",
    67 => x"055334ad",
    68 => x"8408ff05",
    69 => x"ad840cad",
    70 => x"84088025",
    71 => x"eb38ad80",
    72 => x"08ff05ad",
    73 => x"800cad80",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bad80",
    94 => x"08258f38",
    95 => x"82b22dad",
    96 => x"8008ff05",
    97 => x"ad800c82",
    98 => x"f404ad80",
    99 => x"08ad8408",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38ad8008",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134ad",
   108 => x"84088105",
   109 => x"ad840cad",
   110 => x"8408519f",
   111 => x"7125e238",
   112 => x"800bad84",
   113 => x"0cad8008",
   114 => x"8105ad80",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"ad840881",
   120 => x"05ad840c",
   121 => x"ad8408a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"ad840cad",
   125 => x"80088105",
   126 => x"ad800c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bad",
   155 => x"880cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bad88",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"ad880884",
   167 => x"07ad880c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0bab",
   172 => x"bc0c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cad8808",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f8050d",
   198 => x"b1fc0882",
   199 => x"06abe00b",
   200 => x"80f52d52",
   201 => x"5270802e",
   202 => x"85387181",
   203 => x"0752abec",
   204 => x"0b80f52d",
   205 => x"5170802e",
   206 => x"85387184",
   207 => x"075271ac",
   208 => x"f00c0288",
   209 => x"050d0402",
   210 => x"f4050d74",
   211 => x"708206b1",
   212 => x"fc0cabd8",
   213 => x"71810654",
   214 => x"54517188",
   215 => x"1481b72d",
   216 => x"70822a70",
   217 => x"81065151",
   218 => x"70941481",
   219 => x"b72d70ac",
   220 => x"f00c028c",
   221 => x"050d0402",
   222 => x"d4050d7c",
   223 => x"a9c05255",
   224 => x"85f32d99",
   225 => x"d72dacf0",
   226 => x"08802e82",
   227 => x"ca388694",
   228 => x"2dacf008",
   229 => x"538ca72d",
   230 => x"acf00854",
   231 => x"acf00880",
   232 => x"2e82b638",
   233 => x"840bfec4",
   234 => x"0ca9d852",
   235 => x"ad905192",
   236 => x"b92dacf0",
   237 => x"08802e80",
   238 => x"ca387482",
   239 => x"2e098106",
   240 => x"a63872ad",
   241 => x"9c0cada0",
   242 => x"5480fd53",
   243 => x"80747084",
   244 => x"05560cff",
   245 => x"13537280",
   246 => x"25f238ad",
   247 => x"9c52ad90",
   248 => x"5195a42d",
   249 => x"88830474",
   250 => x"812e0981",
   251 => x"069538ad",
   252 => x"9c52ad90",
   253 => x"5194fe2d",
   254 => x"ad9c0870",
   255 => x"fec00c51",
   256 => x"86c72da9",
   257 => x"e452ad90",
   258 => x"5192b92d",
   259 => x"acf00880",
   260 => x"2e81c438",
   261 => x"a9f05185",
   262 => x"f32dad94",
   263 => x"08578077",
   264 => x"595a767a",
   265 => x"2e8b3881",
   266 => x"1a78812a",
   267 => x"595a77f7",
   268 => x"38f71a77",
   269 => x"9fff0654",
   270 => x"5a72802e",
   271 => x"8b38fc80",
   272 => x"17ad9052",
   273 => x"5794d12d",
   274 => x"80772581",
   275 => x"80387952",
   276 => x"77518480",
   277 => x"2dad9c52",
   278 => x"ad905194",
   279 => x"fe2dacf0",
   280 => x"0853acf0",
   281 => x"08802e80",
   282 => x"c938ad9c",
   283 => x"5b805989",
   284 => x"9f047a70",
   285 => x"84055c08",
   286 => x"7081ff06",
   287 => x"71882c70",
   288 => x"81ff0673",
   289 => x"902c7081",
   290 => x"ff067598",
   291 => x"2afec80c",
   292 => x"fec80c58",
   293 => x"fec80c57",
   294 => x"fec80c84",
   295 => x"1a5a5376",
   296 => x"53848077",
   297 => x"25843884",
   298 => x"80537279",
   299 => x"24c43889",
   300 => x"bd04aa80",
   301 => x"5185f32d",
   302 => x"725489d9",
   303 => x"04ad9051",
   304 => x"94d12dfc",
   305 => x"80178119",
   306 => x"595788c8",
   307 => x"04820bfe",
   308 => x"c40c8154",
   309 => x"89d90480",
   310 => x"5473acf0",
   311 => x"0c02ac05",
   312 => x"0d0402f8",
   313 => x"050da1fa",
   314 => x"2d81f72d",
   315 => x"815184e5",
   316 => x"2dfec452",
   317 => x"81720c9f",
   318 => x"c02d9fc0",
   319 => x"2d84720c",
   320 => x"735186f7",
   321 => x"2dabc051",
   322 => x"a3d82d80",
   323 => x"5184e52d",
   324 => x"0288050d",
   325 => x"0402fc05",
   326 => x"0d825189",
   327 => x"e22d0284",
   328 => x"050d0402",
   329 => x"fc050d80",
   330 => x"5189e22d",
   331 => x"0284050d",
   332 => x"0402f405",
   333 => x"0d805186",
   334 => x"c72d810b",
   335 => x"fec40c80",
   336 => x"0bfec00c",
   337 => x"840bfec4",
   338 => x"0c830bfe",
   339 => x"cc0c9fdb",
   340 => x"2da1ee2d",
   341 => x"9fc02d9f",
   342 => x"c02d81f7",
   343 => x"2d815184",
   344 => x"e52d9fc0",
   345 => x"2d9fc02d",
   346 => x"815184e5",
   347 => x"2d815186",
   348 => x"f72dacf0",
   349 => x"08802e80",
   350 => x"db388051",
   351 => x"84e52dab",
   352 => x"c051a3d8",
   353 => x"2d9ff32d",
   354 => x"a3e82dac",
   355 => x"f0085386",
   356 => x"942dacf0",
   357 => x"08fec00c",
   358 => x"86942dac",
   359 => x"f008ad8c",
   360 => x"082e9c38",
   361 => x"acf008ad",
   362 => x"8c0c8452",
   363 => x"725184e5",
   364 => x"2d9fc02d",
   365 => x"9fc02dff",
   366 => x"12527180",
   367 => x"25ee3872",
   368 => x"802e8938",
   369 => x"8a0bfec4",
   370 => x"0c8b8504",
   371 => x"820bfec4",
   372 => x"0c8b8504",
   373 => x"aa905185",
   374 => x"f32d820b",
   375 => x"fec40c80",
   376 => x"0bacf00c",
   377 => x"028c050d",
   378 => x"0402e805",
   379 => x"0d77797b",
   380 => x"58555580",
   381 => x"53727625",
   382 => x"a3387470",
   383 => x"81055680",
   384 => x"f52d7470",
   385 => x"81055680",
   386 => x"f52d5252",
   387 => x"71712e86",
   388 => x"3881518c",
   389 => x"9e048113",
   390 => x"538bf504",
   391 => x"805170ac",
   392 => x"f00c0298",
   393 => x"050d0402",
   394 => x"d8050d80",
   395 => x"0bb1a40c",
   396 => x"ad9c5280",
   397 => x"519cbf2d",
   398 => x"acf00854",
   399 => x"acf0088c",
   400 => x"38aaa851",
   401 => x"85f32d73",
   402 => x"5591c204",
   403 => x"8056810b",
   404 => x"b1c80c88",
   405 => x"53aab452",
   406 => x"add2518b",
   407 => x"e92dacf0",
   408 => x"08762e09",
   409 => x"81068738",
   410 => x"acf008b1",
   411 => x"c80c8853",
   412 => x"aac052ad",
   413 => x"ee518be9",
   414 => x"2dacf008",
   415 => x"8738acf0",
   416 => x"08b1c80c",
   417 => x"b1c80880",
   418 => x"2e80f638",
   419 => x"b0e20b80",
   420 => x"f52db0e3",
   421 => x"0b80f52d",
   422 => x"71982b71",
   423 => x"902b07b0",
   424 => x"e40b80f5",
   425 => x"2d70882b",
   426 => x"7207b0e5",
   427 => x"0b80f52d",
   428 => x"7107b19a",
   429 => x"0b80f52d",
   430 => x"b19b0b80",
   431 => x"f52d7188",
   432 => x"2b07535f",
   433 => x"54525a56",
   434 => x"57557381",
   435 => x"abaa2e09",
   436 => x"81068d38",
   437 => x"75519dda",
   438 => x"2dacf008",
   439 => x"568ded04",
   440 => x"7382d4d5",
   441 => x"2e8738aa",
   442 => x"cc518eae",
   443 => x"04ad9c52",
   444 => x"75519cbf",
   445 => x"2dacf008",
   446 => x"55acf008",
   447 => x"802e83c2",
   448 => x"388853aa",
   449 => x"c052adee",
   450 => x"518be92d",
   451 => x"acf00889",
   452 => x"38810bb1",
   453 => x"a40c8eb4",
   454 => x"048853aa",
   455 => x"b452add2",
   456 => x"518be92d",
   457 => x"acf00880",
   458 => x"2e8a38aa",
   459 => x"e05185f3",
   460 => x"2d8f8e04",
   461 => x"b19a0b80",
   462 => x"f52d5473",
   463 => x"80d52e09",
   464 => x"810680ca",
   465 => x"38b19b0b",
   466 => x"80f52d54",
   467 => x"7381aa2e",
   468 => x"098106ba",
   469 => x"38800bad",
   470 => x"9c0b80f5",
   471 => x"2d565474",
   472 => x"81e92e83",
   473 => x"38815474",
   474 => x"81eb2e8c",
   475 => x"38805573",
   476 => x"752e0981",
   477 => x"0682cb38",
   478 => x"ada70b80",
   479 => x"f52d5574",
   480 => x"8d38ada8",
   481 => x"0b80f52d",
   482 => x"5473822e",
   483 => x"86388055",
   484 => x"91c204ad",
   485 => x"a90b80f5",
   486 => x"2d70b19c",
   487 => x"0cff05b1",
   488 => x"a00cadaa",
   489 => x"0b80f52d",
   490 => x"adab0b80",
   491 => x"f52d5876",
   492 => x"05778280",
   493 => x"290570b1",
   494 => x"a80cadac",
   495 => x"0b80f52d",
   496 => x"70b1bc0c",
   497 => x"b1a40859",
   498 => x"57587680",
   499 => x"2e81a338",
   500 => x"8853aac0",
   501 => x"52adee51",
   502 => x"8be92dac",
   503 => x"f00881e2",
   504 => x"38b19c08",
   505 => x"70842bb1",
   506 => x"c00c70b1",
   507 => x"b80cadc1",
   508 => x"0b80f52d",
   509 => x"adc00b80",
   510 => x"f52d7182",
   511 => x"802905ad",
   512 => x"c20b80f5",
   513 => x"2d708480",
   514 => x"802912ad",
   515 => x"c30b80f5",
   516 => x"2d708180",
   517 => x"0a291270",
   518 => x"b1c40cb1",
   519 => x"bc087129",
   520 => x"b1a80805",
   521 => x"70b1ac0c",
   522 => x"adc90b80",
   523 => x"f52dadc8",
   524 => x"0b80f52d",
   525 => x"71828029",
   526 => x"05adca0b",
   527 => x"80f52d70",
   528 => x"84808029",
   529 => x"12adcb0b",
   530 => x"80f52d70",
   531 => x"982b81f0",
   532 => x"0a067205",
   533 => x"70b1b00c",
   534 => x"fe117e29",
   535 => x"7705b1b4",
   536 => x"0c525952",
   537 => x"43545e51",
   538 => x"5259525d",
   539 => x"57595791",
   540 => x"c004adae",
   541 => x"0b80f52d",
   542 => x"adad0b80",
   543 => x"f52d7182",
   544 => x"80290570",
   545 => x"b1c00c70",
   546 => x"a02983ff",
   547 => x"0570892a",
   548 => x"70b1b80c",
   549 => x"adb30b80",
   550 => x"f52dadb2",
   551 => x"0b80f52d",
   552 => x"71828029",
   553 => x"0570b1c4",
   554 => x"0c7b7129",
   555 => x"1e70b1b4",
   556 => x"0c7db1b0",
   557 => x"0c7305b1",
   558 => x"ac0c555e",
   559 => x"51515555",
   560 => x"815574ac",
   561 => x"f00c02a8",
   562 => x"050d0402",
   563 => x"ec050d76",
   564 => x"70872c71",
   565 => x"80ff0655",
   566 => x"5654b1a4",
   567 => x"088a3873",
   568 => x"882c7481",
   569 => x"ff065455",
   570 => x"ad9c52b1",
   571 => x"a8081551",
   572 => x"9cbf2dac",
   573 => x"f00854ac",
   574 => x"f008802e",
   575 => x"b338b1a4",
   576 => x"08802e98",
   577 => x"38728429",
   578 => x"ad9c0570",
   579 => x"0852539d",
   580 => x"da2dacf0",
   581 => x"08f00a06",
   582 => x"5392ae04",
   583 => x"7210ad9c",
   584 => x"057080e0",
   585 => x"2d52539e",
   586 => x"8a2dacf0",
   587 => x"08537254",
   588 => x"73acf00c",
   589 => x"0294050d",
   590 => x"0402c805",
   591 => x"0d7f615f",
   592 => x"5b800bb1",
   593 => x"b008b1b4",
   594 => x"08595d56",
   595 => x"b1a40876",
   596 => x"2e8a38b1",
   597 => x"9c08842b",
   598 => x"5892e204",
   599 => x"b1b80884",
   600 => x"2b588059",
   601 => x"78782781",
   602 => x"a938788f",
   603 => x"06a01757",
   604 => x"54738f38",
   605 => x"ad9c5276",
   606 => x"51811757",
   607 => x"9cbf2dad",
   608 => x"9c568076",
   609 => x"80f52d56",
   610 => x"5474742e",
   611 => x"83388154",
   612 => x"7481e52e",
   613 => x"80f63881",
   614 => x"70750655",
   615 => x"5d73802e",
   616 => x"80ea388b",
   617 => x"1680f52d",
   618 => x"98065a79",
   619 => x"80de388b",
   620 => x"537d5275",
   621 => x"518be92d",
   622 => x"acf00880",
   623 => x"cf389c16",
   624 => x"08519dda",
   625 => x"2dacf008",
   626 => x"841c0c9a",
   627 => x"1680e02d",
   628 => x"519e8a2d",
   629 => x"acf008ac",
   630 => x"f008881d",
   631 => x"0cacf008",
   632 => x"5555b1a4",
   633 => x"08802e98",
   634 => x"38941680",
   635 => x"e02d519e",
   636 => x"8a2dacf0",
   637 => x"08902b83",
   638 => x"fff00a06",
   639 => x"70165154",
   640 => x"73881c0c",
   641 => x"797b0c7c",
   642 => x"5494c804",
   643 => x"81195992",
   644 => x"e404b1a4",
   645 => x"08802eae",
   646 => x"387b5191",
   647 => x"cb2dacf0",
   648 => x"08acf008",
   649 => x"80ffffff",
   650 => x"f806555c",
   651 => x"7380ffff",
   652 => x"fff82e92",
   653 => x"38acf008",
   654 => x"fe05b19c",
   655 => x"0829b1ac",
   656 => x"08055792",
   657 => x"e2048054",
   658 => x"73acf00c",
   659 => x"02b8050d",
   660 => x"0402f405",
   661 => x"0d747008",
   662 => x"8105710c",
   663 => x"7008b1a0",
   664 => x"08065353",
   665 => x"718e3888",
   666 => x"13085191",
   667 => x"cb2dacf0",
   668 => x"0888140c",
   669 => x"810bacf0",
   670 => x"0c028c05",
   671 => x"0d0402f0",
   672 => x"050d7588",
   673 => x"1108fe05",
   674 => x"b19c0829",
   675 => x"b1ac0811",
   676 => x"7208b1a0",
   677 => x"08060579",
   678 => x"55535454",
   679 => x"9cbf2d02",
   680 => x"90050d04",
   681 => x"02f0050d",
   682 => x"75881108",
   683 => x"fe05b19c",
   684 => x"0829b1ac",
   685 => x"08117208",
   686 => x"b1a00806",
   687 => x"05795553",
   688 => x"54549aff",
   689 => x"2d029005",
   690 => x"0d0402f4",
   691 => x"050dd452",
   692 => x"81ff720c",
   693 => x"71085381",
   694 => x"ff720c72",
   695 => x"882b83fe",
   696 => x"80067208",
   697 => x"7081ff06",
   698 => x"51525381",
   699 => x"ff720c72",
   700 => x"7107882b",
   701 => x"72087081",
   702 => x"ff065152",
   703 => x"5381ff72",
   704 => x"0c727107",
   705 => x"882b7208",
   706 => x"7081ff06",
   707 => x"7207acf0",
   708 => x"0c525302",
   709 => x"8c050d04",
   710 => x"02f4050d",
   711 => x"74767181",
   712 => x"ff06d40c",
   713 => x"5353b1cc",
   714 => x"08853871",
   715 => x"892b5271",
   716 => x"982ad40c",
   717 => x"71902a70",
   718 => x"81ff06d4",
   719 => x"0c517188",
   720 => x"2a7081ff",
   721 => x"06d40c51",
   722 => x"7181ff06",
   723 => x"d40c7290",
   724 => x"2a7081ff",
   725 => x"06d40c51",
   726 => x"d4087081",
   727 => x"ff065151",
   728 => x"82b8bf52",
   729 => x"7081ff2e",
   730 => x"09810694",
   731 => x"3881ff0b",
   732 => x"d40cd408",
   733 => x"7081ff06",
   734 => x"ff145451",
   735 => x"5171e538",
   736 => x"70acf00c",
   737 => x"028c050d",
   738 => x"0402fc05",
   739 => x"0d81c751",
   740 => x"81ff0bd4",
   741 => x"0cff1151",
   742 => x"708025f4",
   743 => x"38028405",
   744 => x"0d0402f0",
   745 => x"050d9789",
   746 => x"2d8fcf53",
   747 => x"805287fc",
   748 => x"80f75196",
   749 => x"982dacf0",
   750 => x"0854acf0",
   751 => x"08812e09",
   752 => x"8106a338",
   753 => x"81ff0bd4",
   754 => x"0c820a52",
   755 => x"849c80e9",
   756 => x"5196982d",
   757 => x"acf0088b",
   758 => x"3881ff0b",
   759 => x"d40c7353",
   760 => x"97ec0497",
   761 => x"892dff13",
   762 => x"5372c138",
   763 => x"72acf00c",
   764 => x"0290050d",
   765 => x"0402f405",
   766 => x"0d81ff0b",
   767 => x"d40c9353",
   768 => x"805287fc",
   769 => x"80c15196",
   770 => x"982dacf0",
   771 => x"088b3881",
   772 => x"ff0bd40c",
   773 => x"815398a2",
   774 => x"0497892d",
   775 => x"ff135372",
   776 => x"df3872ac",
   777 => x"f00c028c",
   778 => x"050d0402",
   779 => x"f0050d97",
   780 => x"892d83aa",
   781 => x"52849c80",
   782 => x"c8519698",
   783 => x"2dacf008",
   784 => x"812e0981",
   785 => x"06923895",
   786 => x"ca2dacf0",
   787 => x"0883ffff",
   788 => x"06537283",
   789 => x"aa2e9738",
   790 => x"97f52d98",
   791 => x"e9048154",
   792 => x"99ce04aa",
   793 => x"ec5185f3",
   794 => x"2d805499",
   795 => x"ce0481ff",
   796 => x"0bd40cb1",
   797 => x"5397a22d",
   798 => x"acf00880",
   799 => x"2e80c038",
   800 => x"805287fc",
   801 => x"80fa5196",
   802 => x"982dacf0",
   803 => x"08b13881",
   804 => x"ff0bd40c",
   805 => x"d4085381",
   806 => x"ff0bd40c",
   807 => x"81ff0bd4",
   808 => x"0c81ff0b",
   809 => x"d40c81ff",
   810 => x"0bd40c72",
   811 => x"862a7081",
   812 => x"06acf008",
   813 => x"56515372",
   814 => x"802e9338",
   815 => x"98de0472",
   816 => x"822eff9f",
   817 => x"38ff1353",
   818 => x"72ffaa38",
   819 => x"725473ac",
   820 => x"f00c0290",
   821 => x"050d0402",
   822 => x"f0050d81",
   823 => x"0bb1cc0c",
   824 => x"8454d008",
   825 => x"708f2a70",
   826 => x"81065151",
   827 => x"5372f338",
   828 => x"72d00c97",
   829 => x"892daafc",
   830 => x"5185f32d",
   831 => x"d008708f",
   832 => x"2a708106",
   833 => x"51515372",
   834 => x"f338810b",
   835 => x"d00cb153",
   836 => x"805284d4",
   837 => x"80c05196",
   838 => x"982dacf0",
   839 => x"08812ea1",
   840 => x"3872822e",
   841 => x"0981068c",
   842 => x"38ab8851",
   843 => x"85f32d80",
   844 => x"539af604",
   845 => x"ff135372",
   846 => x"d738ff14",
   847 => x"5473ffa2",
   848 => x"3898ab2d",
   849 => x"acf008b1",
   850 => x"cc0cacf0",
   851 => x"088b3881",
   852 => x"5287fc80",
   853 => x"d0519698",
   854 => x"2d81ff0b",
   855 => x"d40cd008",
   856 => x"708f2a70",
   857 => x"81065151",
   858 => x"5372f338",
   859 => x"72d00c81",
   860 => x"ff0bd40c",
   861 => x"815372ac",
   862 => x"f00c0290",
   863 => x"050d0402",
   864 => x"e8050d78",
   865 => x"5681ff0b",
   866 => x"d40cd008",
   867 => x"708f2a70",
   868 => x"81065151",
   869 => x"5372f338",
   870 => x"82810bd0",
   871 => x"0c81ff0b",
   872 => x"d40c7752",
   873 => x"87fc80d8",
   874 => x"5196982d",
   875 => x"acf00880",
   876 => x"2e8c38ab",
   877 => x"a05185f3",
   878 => x"2d81539c",
   879 => x"b60481ff",
   880 => x"0bd40c81",
   881 => x"fe0bd40c",
   882 => x"80ff5575",
   883 => x"70840557",
   884 => x"0870982a",
   885 => x"d40c7090",
   886 => x"2c7081ff",
   887 => x"06d40c54",
   888 => x"70882c70",
   889 => x"81ff06d4",
   890 => x"0c547081",
   891 => x"ff06d40c",
   892 => x"54ff1555",
   893 => x"748025d3",
   894 => x"3881ff0b",
   895 => x"d40c81ff",
   896 => x"0bd40c81",
   897 => x"ff0bd40c",
   898 => x"868da054",
   899 => x"81ff0bd4",
   900 => x"0cd40881",
   901 => x"ff065574",
   902 => x"8738ff14",
   903 => x"5473ed38",
   904 => x"81ff0bd4",
   905 => x"0cd00870",
   906 => x"8f2a7081",
   907 => x"06515153",
   908 => x"72f33872",
   909 => x"d00c72ac",
   910 => x"f00c0298",
   911 => x"050d0402",
   912 => x"e8050d78",
   913 => x"55805681",
   914 => x"ff0bd40c",
   915 => x"d008708f",
   916 => x"2a708106",
   917 => x"51515372",
   918 => x"f3388281",
   919 => x"0bd00c81",
   920 => x"ff0bd40c",
   921 => x"775287fc",
   922 => x"80d15196",
   923 => x"982d80db",
   924 => x"c6df54ac",
   925 => x"f008802e",
   926 => x"8a38aa80",
   927 => x"5185f32d",
   928 => x"9dd10481",
   929 => x"ff0bd40c",
   930 => x"d4087081",
   931 => x"ff065153",
   932 => x"7281fe2e",
   933 => x"0981069d",
   934 => x"3880ff53",
   935 => x"95ca2dac",
   936 => x"f0087570",
   937 => x"8405570c",
   938 => x"ff135372",
   939 => x"8025ed38",
   940 => x"81569dbb",
   941 => x"04ff1454",
   942 => x"73c93881",
   943 => x"ff0bd40c",
   944 => x"d008708f",
   945 => x"2a708106",
   946 => x"51515372",
   947 => x"f33872d0",
   948 => x"0c75acf0",
   949 => x"0c029805",
   950 => x"0d0402f4",
   951 => x"050d7470",
   952 => x"882a83fe",
   953 => x"80067072",
   954 => x"982a0772",
   955 => x"882b87fc",
   956 => x"80800673",
   957 => x"982b81f0",
   958 => x"0a067173",
   959 => x"0707acf0",
   960 => x"0c565153",
   961 => x"51028c05",
   962 => x"0d0402f8",
   963 => x"050d028e",
   964 => x"0580f52d",
   965 => x"74882b07",
   966 => x"7083ffff",
   967 => x"06acf00c",
   968 => x"51028805",
   969 => x"0d0402fc",
   970 => x"050d7251",
   971 => x"80710c80",
   972 => x"0b84120c",
   973 => x"0284050d",
   974 => x"0402f005",
   975 => x"0d757008",
   976 => x"84120853",
   977 => x"5353ff54",
   978 => x"71712ea8",
   979 => x"38a1f42d",
   980 => x"84130870",
   981 => x"84291488",
   982 => x"11700870",
   983 => x"81ff0684",
   984 => x"18088111",
   985 => x"8706841a",
   986 => x"0c535155",
   987 => x"515151a1",
   988 => x"ee2d7154",
   989 => x"73acf00c",
   990 => x"0290050d",
   991 => x"0402f805",
   992 => x"0da1f42d",
   993 => x"e008708b",
   994 => x"2a708106",
   995 => x"51525270",
   996 => x"802e9d38",
   997 => x"b1d00870",
   998 => x"8429b1d8",
   999 => x"057381ff",
  1000 => x"06710c51",
  1001 => x"51b1d008",
  1002 => x"81118706",
  1003 => x"b1d00c51",
  1004 => x"800bb1f8",
  1005 => x"0ca1e72d",
  1006 => x"a1ee2d02",
  1007 => x"88050d04",
  1008 => x"02fc050d",
  1009 => x"a1f42d81",
  1010 => x"0bb1f80c",
  1011 => x"a1ee2db1",
  1012 => x"f8085170",
  1013 => x"fa380284",
  1014 => x"050d0402",
  1015 => x"fc050db1",
  1016 => x"d0519ea6",
  1017 => x"2d9efd51",
  1018 => x"a1e32da1",
  1019 => x"8d2d0284",
  1020 => x"050d0402",
  1021 => x"f4050da0",
  1022 => x"f504acf0",
  1023 => x"0881f02e",
  1024 => x"09810689",
  1025 => x"38810bac",
  1026 => x"e40ca0f5",
  1027 => x"04acf008",
  1028 => x"81e02e09",
  1029 => x"81068938",
  1030 => x"810bace8",
  1031 => x"0ca0f504",
  1032 => x"acf00852",
  1033 => x"ace80880",
  1034 => x"2e8838ac",
  1035 => x"f0088180",
  1036 => x"05527184",
  1037 => x"2c728f06",
  1038 => x"5353ace4",
  1039 => x"08802e99",
  1040 => x"38728429",
  1041 => x"aca40572",
  1042 => x"1381712b",
  1043 => x"70097308",
  1044 => x"06730c51",
  1045 => x"5353a0eb",
  1046 => x"04728429",
  1047 => x"aca40572",
  1048 => x"1383712b",
  1049 => x"72080772",
  1050 => x"0c535380",
  1051 => x"0bace80c",
  1052 => x"800bace4",
  1053 => x"0cb1d051",
  1054 => x"9eb92dac",
  1055 => x"f008ff24",
  1056 => x"fef83880",
  1057 => x"0bacf00c",
  1058 => x"028c050d",
  1059 => x"0402f805",
  1060 => x"0daca452",
  1061 => x"8f518072",
  1062 => x"70840554",
  1063 => x"0cff1151",
  1064 => x"708025f2",
  1065 => x"38028805",
  1066 => x"0d0402f0",
  1067 => x"050d7551",
  1068 => x"a1f42d70",
  1069 => x"822cfc06",
  1070 => x"aca41172",
  1071 => x"109e0671",
  1072 => x"0870722a",
  1073 => x"70830682",
  1074 => x"742b7009",
  1075 => x"7406760c",
  1076 => x"54515657",
  1077 => x"535153a1",
  1078 => x"ee2d71ac",
  1079 => x"f00c0290",
  1080 => x"050d0471",
  1081 => x"980c04ff",
  1082 => x"b008acf0",
  1083 => x"0c04810b",
  1084 => x"ffb00c04",
  1085 => x"800bffb0",
  1086 => x"0c0402fc",
  1087 => x"050d800b",
  1088 => x"acec0c80",
  1089 => x"5184e52d",
  1090 => x"0284050d",
  1091 => x"0402ec05",
  1092 => x"0d765480",
  1093 => x"52870b88",
  1094 => x"1580f52d",
  1095 => x"56537472",
  1096 => x"248338a0",
  1097 => x"53725182",
  1098 => x"ee2d8112",
  1099 => x"8b1580f5",
  1100 => x"2d545272",
  1101 => x"7225de38",
  1102 => x"0294050d",
  1103 => x"0402f005",
  1104 => x"0db28008",
  1105 => x"5481f72d",
  1106 => x"800bb284",
  1107 => x"0c730880",
  1108 => x"2e818038",
  1109 => x"820bad84",
  1110 => x"0cb28408",
  1111 => x"8f06ad80",
  1112 => x"0c730852",
  1113 => x"71832e96",
  1114 => x"38718326",
  1115 => x"89387181",
  1116 => x"2eaf38a3",
  1117 => x"be047185",
  1118 => x"2e9f38a3",
  1119 => x"be048814",
  1120 => x"80f52d84",
  1121 => x"1508abb0",
  1122 => x"53545285",
  1123 => x"f32d7184",
  1124 => x"29137008",
  1125 => x"5252a3c2",
  1126 => x"047351a2",
  1127 => x"8d2da3be",
  1128 => x"04b1fc08",
  1129 => x"8815082c",
  1130 => x"70810651",
  1131 => x"5271802e",
  1132 => x"8738abb4",
  1133 => x"51a3bb04",
  1134 => x"abb85185",
  1135 => x"f32d8414",
  1136 => x"085185f3",
  1137 => x"2db28408",
  1138 => x"8105b284",
  1139 => x"0c8c1454",
  1140 => x"a2cd0402",
  1141 => x"90050d04",
  1142 => x"71b2800c",
  1143 => x"a2bd2db2",
  1144 => x"8408ff05",
  1145 => x"b2880c04",
  1146 => x"02ec050d",
  1147 => x"b2800855",
  1148 => x"80f851a1",
  1149 => x"aa2dacf0",
  1150 => x"08812a70",
  1151 => x"81065152",
  1152 => x"719b3887",
  1153 => x"51a1aa2d",
  1154 => x"acf00881",
  1155 => x"2a708106",
  1156 => x"51527180",
  1157 => x"2eb138a4",
  1158 => x"9d049ff3",
  1159 => x"2d8751a1",
  1160 => x"aa2dacf0",
  1161 => x"08f438a4",
  1162 => x"ad049ff3",
  1163 => x"2d80f851",
  1164 => x"a1aa2dac",
  1165 => x"f008f338",
  1166 => x"acec0881",
  1167 => x"3270acec",
  1168 => x"0c705252",
  1169 => x"84e52dac",
  1170 => x"ec08a238",
  1171 => x"80da51a1",
  1172 => x"aa2d81f5",
  1173 => x"51a1aa2d",
  1174 => x"81f251a1",
  1175 => x"aa2d81eb",
  1176 => x"51a1aa2d",
  1177 => x"81f451a1",
  1178 => x"aa2da8b1",
  1179 => x"0481f551",
  1180 => x"a1aa2dac",
  1181 => x"f008812a",
  1182 => x"70810651",
  1183 => x"5271802e",
  1184 => x"8f38b288",
  1185 => x"08527180",
  1186 => x"2e8638ff",
  1187 => x"12b2880c",
  1188 => x"81f251a1",
  1189 => x"aa2dacf0",
  1190 => x"08812a70",
  1191 => x"81065152",
  1192 => x"71802e95",
  1193 => x"38b28408",
  1194 => x"ff05b288",
  1195 => x"08545272",
  1196 => x"72258638",
  1197 => x"8113b288",
  1198 => x"0cb28808",
  1199 => x"70535473",
  1200 => x"802e8a38",
  1201 => x"8c15ff15",
  1202 => x"5555a5bf",
  1203 => x"04820bad",
  1204 => x"840c718f",
  1205 => x"06ad800c",
  1206 => x"81eb51a1",
  1207 => x"aa2dacf0",
  1208 => x"08812a70",
  1209 => x"81065152",
  1210 => x"71802ead",
  1211 => x"38740885",
  1212 => x"2e098106",
  1213 => x"a4388815",
  1214 => x"80f52dff",
  1215 => x"05527188",
  1216 => x"1681b72d",
  1217 => x"71982b52",
  1218 => x"71802588",
  1219 => x"38800b88",
  1220 => x"1681b72d",
  1221 => x"7451a28d",
  1222 => x"2d81f451",
  1223 => x"a1aa2dac",
  1224 => x"f008812a",
  1225 => x"70810651",
  1226 => x"5271802e",
  1227 => x"b3387408",
  1228 => x"852e0981",
  1229 => x"06aa3888",
  1230 => x"1580f52d",
  1231 => x"81055271",
  1232 => x"881681b7",
  1233 => x"2d7181ff",
  1234 => x"068b1680",
  1235 => x"f52d5452",
  1236 => x"72722787",
  1237 => x"38728816",
  1238 => x"81b72d74",
  1239 => x"51a28d2d",
  1240 => x"80da51a1",
  1241 => x"aa2dacf0",
  1242 => x"08812a70",
  1243 => x"81065152",
  1244 => x"71802e80",
  1245 => x"fb38b280",
  1246 => x"08b28808",
  1247 => x"55537380",
  1248 => x"2e8a388c",
  1249 => x"13ff1555",
  1250 => x"53a6fe04",
  1251 => x"72085271",
  1252 => x"822ea638",
  1253 => x"71822689",
  1254 => x"3871812e",
  1255 => x"a538a7f0",
  1256 => x"0471832e",
  1257 => x"ad387184",
  1258 => x"2e098106",
  1259 => x"80c23888",
  1260 => x"130851a3",
  1261 => x"d82da7f0",
  1262 => x"04881308",
  1263 => x"52712da7",
  1264 => x"f004810b",
  1265 => x"8814082b",
  1266 => x"b1fc0832",
  1267 => x"b1fc0ca7",
  1268 => x"ed048813",
  1269 => x"80f52d81",
  1270 => x"058b1480",
  1271 => x"f52d5354",
  1272 => x"71742483",
  1273 => x"38805473",
  1274 => x"881481b7",
  1275 => x"2da2bd2d",
  1276 => x"8054800b",
  1277 => x"ad840c73",
  1278 => x"8f06ad80",
  1279 => x"0ca05273",
  1280 => x"b288082e",
  1281 => x"09810698",
  1282 => x"38b28408",
  1283 => x"ff057432",
  1284 => x"70098105",
  1285 => x"7072079f",
  1286 => x"2a917131",
  1287 => x"51515353",
  1288 => x"715182ee",
  1289 => x"2d811454",
  1290 => x"8e7425c6",
  1291 => x"38acec08",
  1292 => x"5271acf0",
  1293 => x"0c029405",
  1294 => x"0d040000",
  1295 => x"00ffffff",
  1296 => x"ff00ffff",
  1297 => x"ffff00ff",
  1298 => x"ffffff00",
  1299 => x"52657365",
  1300 => x"74000000",
  1301 => x"53617665",
  1302 => x"20616e64",
  1303 => x"20526573",
  1304 => x"65740000",
  1305 => x"5363616e",
  1306 => x"6c696e65",
  1307 => x"73000000",
  1308 => x"45786974",
  1309 => x"00000000",
  1310 => x"50432045",
  1311 => x"6e67696e",
  1312 => x"65206d6f",
  1313 => x"64650000",
  1314 => x"54757262",
  1315 => x"6f677261",
  1316 => x"66782031",
  1317 => x"36206d6f",
  1318 => x"64650000",
  1319 => x"56474120",
  1320 => x"2d203331",
  1321 => x"4b487a2c",
  1322 => x"20363048",
  1323 => x"7a000000",
  1324 => x"5456202d",
  1325 => x"20343830",
  1326 => x"692c2036",
  1327 => x"30487a00",
  1328 => x"496e6974",
  1329 => x"69616c69",
  1330 => x"7a696e67",
  1331 => x"20534420",
  1332 => x"63617264",
  1333 => x"0a000000",
  1334 => x"46504741",
  1335 => x"50434520",
  1336 => x"43464700",
  1337 => x"4d535833",
  1338 => x"42494f53",
  1339 => x"53595300",
  1340 => x"4c6f6164",
  1341 => x"696e6720",
  1342 => x"524f4d0a",
  1343 => x"00000000",
  1344 => x"52656164",
  1345 => x"20666169",
  1346 => x"6c65640a",
  1347 => x"00000000",
  1348 => x"4c6f6164",
  1349 => x"696e6720",
  1350 => x"42494f53",
  1351 => x"20666169",
  1352 => x"6c65640a",
  1353 => x"00000000",
  1354 => x"4d425220",
  1355 => x"6661696c",
  1356 => x"0a000000",
  1357 => x"46415431",
  1358 => x"36202020",
  1359 => x"00000000",
  1360 => x"46415433",
  1361 => x"32202020",
  1362 => x"00000000",
  1363 => x"4e6f2070",
  1364 => x"61727469",
  1365 => x"74696f6e",
  1366 => x"20736967",
  1367 => x"0a000000",
  1368 => x"42616420",
  1369 => x"70617274",
  1370 => x"0a000000",
  1371 => x"53444843",
  1372 => x"20657272",
  1373 => x"6f72210a",
  1374 => x"00000000",
  1375 => x"53442069",
  1376 => x"6e69742e",
  1377 => x"2e2e0a00",
  1378 => x"53442063",
  1379 => x"61726420",
  1380 => x"72657365",
  1381 => x"74206661",
  1382 => x"696c6564",
  1383 => x"210a0000",
  1384 => x"57726974",
  1385 => x"65206661",
  1386 => x"696c6564",
  1387 => x"0a000000",
  1388 => x"16200000",
  1389 => x"14200000",
  1390 => x"15200000",
  1391 => x"00000002",
  1392 => x"00000002",
  1393 => x"0000144c",
  1394 => x"00000523",
  1395 => x"00000002",
  1396 => x"00001454",
  1397 => x"00000515",
  1398 => x"00000003",
  1399 => x"0000161c",
  1400 => x"00000002",
  1401 => x"00000001",
  1402 => x"00001464",
  1403 => x"00000001",
  1404 => x"00000003",
  1405 => x"00001614",
  1406 => x"00000002",
  1407 => x"00000002",
  1408 => x"00001470",
  1409 => x"000010fa",
  1410 => x"00000000",
  1411 => x"00000000",
  1412 => x"00000000",
  1413 => x"00001478",
  1414 => x"00001488",
  1415 => x"0000149c",
  1416 => x"000014b0",
  1417 => x"00000000",
  1418 => x"00000000",
  1419 => x"00000000",
  1420 => x"00000000",
  1421 => x"00000000",
  1422 => x"00000000",
  1423 => x"00000000",
  1424 => x"00000000",
  1425 => x"00000000",
  1426 => x"00000000",
  1427 => x"00000000",
  1428 => x"00000000",
  1429 => x"00000000",
  1430 => x"00000000",
  1431 => x"00000000",
  1432 => x"00000000",
  1433 => x"00000000",
  1434 => x"00000000",
  1435 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

