-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb5",
     9 => x"b4080b0b",
    10 => x"0bb5b808",
    11 => x"0b0b0bb5",
    12 => x"bc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b5bc0c0b",
    16 => x"0b0bb5b8",
    17 => x"0c0b0b0b",
    18 => x"b5b40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bafa8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b5b470bc",
    57 => x"a8278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8cc50402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b5c40c9f",
    65 => x"0bb5c80c",
    66 => x"a0717081",
    67 => x"055334b5",
    68 => x"c808ff05",
    69 => x"b5c80cb5",
    70 => x"c8088025",
    71 => x"eb38b5c4",
    72 => x"08ff05b5",
    73 => x"c40cb5c4",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb5c4",
    94 => x"08258f38",
    95 => x"82b22db5",
    96 => x"c408ff05",
    97 => x"b5c40c82",
    98 => x"f404b5c4",
    99 => x"08b5c808",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b5c408",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b5",
   108 => x"c8088105",
   109 => x"b5c80cb5",
   110 => x"c808519f",
   111 => x"7125e238",
   112 => x"800bb5c8",
   113 => x"0cb5c408",
   114 => x"8105b5c4",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b5c80881",
   120 => x"05b5c80c",
   121 => x"b5c808a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b5c80cb5",
   125 => x"c4088105",
   126 => x"b5c40c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb5",
   155 => x"cc0cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb5cc",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b5cc0884",
   167 => x"07b5cc0c",
   168 => x"5573842b",
   169 => x"87e87125",
   170 => x"83713170",
   171 => x"0b0b0bb2",
   172 => x"bc0c8171",
   173 => x"2bf6880c",
   174 => x"fea413ff",
   175 => x"122c7888",
   176 => x"29ff9405",
   177 => x"70812cb5",
   178 => x"cc085258",
   179 => x"52555152",
   180 => x"5476802e",
   181 => x"85387081",
   182 => x"075170f6",
   183 => x"940c7109",
   184 => x"8105f680",
   185 => x"0c720981",
   186 => x"05f6840c",
   187 => x"0294050d",
   188 => x"0402f405",
   189 => x"0d745372",
   190 => x"70810554",
   191 => x"80f52d52",
   192 => x"71802e89",
   193 => x"38715182",
   194 => x"ee2d85f7",
   195 => x"04028c05",
   196 => x"0d0402f4",
   197 => x"050d7470",
   198 => x"8206bc90",
   199 => x"0cb2d871",
   200 => x"81065454",
   201 => x"51718814",
   202 => x"81b72d70",
   203 => x"822a7081",
   204 => x"06515170",
   205 => x"941481b7",
   206 => x"2d70b5b4",
   207 => x"0c028c05",
   208 => x"0d0402f4",
   209 => x"050db0c0",
   210 => x"52b5d451",
   211 => x"95de2db5",
   212 => x"b408802e",
   213 => x"9538b7b0",
   214 => x"52b5d451",
   215 => x"98942db7",
   216 => x"b00870fe",
   217 => x"c00c5186",
   218 => x"922d028c",
   219 => x"050d0402",
   220 => x"f8050dbc",
   221 => x"90088206",
   222 => x"b2e00b80",
   223 => x"f52d5252",
   224 => x"70802e85",
   225 => x"38718107",
   226 => x"52b2f80b",
   227 => x"80f52d51",
   228 => x"70802e85",
   229 => x"38718407",
   230 => x"5271b5b4",
   231 => x"0c028805",
   232 => x"0d0402f0",
   233 => x"050d86ef",
   234 => x"2db5b408",
   235 => x"b0c053b5",
   236 => x"d4525395",
   237 => x"de2db5b4",
   238 => x"08802ea3",
   239 => x"3872b7b0",
   240 => x"0cb7b454",
   241 => x"80fd5380",
   242 => x"74708405",
   243 => x"560cff13",
   244 => x"53728025",
   245 => x"f238b7b0",
   246 => x"52b5d451",
   247 => x"98ba2d02",
   248 => x"90050d04",
   249 => x"02d8050d",
   250 => x"810bfec4",
   251 => x"0c840bfe",
   252 => x"c40c7b52",
   253 => x"b5d45195",
   254 => x"de2db5b4",
   255 => x"0853b5b4",
   256 => x"08802e81",
   257 => x"ba38b5d8",
   258 => x"0856800b",
   259 => x"ff175859",
   260 => x"76792e8b",
   261 => x"38811977",
   262 => x"812a5859",
   263 => x"76f738f7",
   264 => x"19769fff",
   265 => x"06545972",
   266 => x"802e8b38",
   267 => x"fc8016b5",
   268 => x"d4525697",
   269 => x"e72d8076",
   270 => x"2580fa38",
   271 => x"78527651",
   272 => x"84802db7",
   273 => x"b052b5d4",
   274 => x"5198942d",
   275 => x"b5b40853",
   276 => x"b5b40880",
   277 => x"2e80c838",
   278 => x"b7b05a80",
   279 => x"58898c04",
   280 => x"79708405",
   281 => x"5b087083",
   282 => x"fe800671",
   283 => x"882b83fe",
   284 => x"80067188",
   285 => x"2a077288",
   286 => x"2a83fe80",
   287 => x"0673982a",
   288 => x"07fec80c",
   289 => x"fec80c56",
   290 => x"84195953",
   291 => x"75538480",
   292 => x"76258438",
   293 => x"84805372",
   294 => x"7824c538",
   295 => x"89a504b0",
   296 => x"cc5189c2",
   297 => x"04b5d451",
   298 => x"97e72dfc",
   299 => x"80168118",
   300 => x"585688b6",
   301 => x"04820bfe",
   302 => x"c40c8153",
   303 => x"89c504b0",
   304 => x"dc5185f1",
   305 => x"2d72b5b4",
   306 => x"0c02a805",
   307 => x"0d0402fc",
   308 => x"050da5a8",
   309 => x"2dfec451",
   310 => x"81710c82",
   311 => x"710c0284",
   312 => x"050d0402",
   313 => x"f4050d74",
   314 => x"10157084",
   315 => x"29b3b405",
   316 => x"70085551",
   317 => x"5272802e",
   318 => x"9b387280",
   319 => x"f52d5271",
   320 => x"802e9138",
   321 => x"b0e45185",
   322 => x"f12d7251",
   323 => x"85f12d72",
   324 => x"5187e42d",
   325 => x"b2c051a7",
   326 => x"862da5a8",
   327 => x"2d805184",
   328 => x"e52d028c",
   329 => x"050d0402",
   330 => x"e8050d80",
   331 => x"70565675",
   332 => x"b4e40825",
   333 => x"af38bbbc",
   334 => x"08762ea8",
   335 => x"38745195",
   336 => x"892db5b4",
   337 => x"08098105",
   338 => x"70b5b408",
   339 => x"079f2a77",
   340 => x"05811757",
   341 => x"575275b4",
   342 => x"e4082588",
   343 => x"38bbbc08",
   344 => x"7526da38",
   345 => x"805674bb",
   346 => x"bc082780",
   347 => x"d0387451",
   348 => x"95892d75",
   349 => x"842b52b5",
   350 => x"b408802e",
   351 => x"ae38b5e0",
   352 => x"128117b5",
   353 => x"b4085657",
   354 => x"528a5373",
   355 => x"70810555",
   356 => x"80f52d72",
   357 => x"70810554",
   358 => x"81b72dff",
   359 => x"13537280",
   360 => x"25e93880",
   361 => x"7281b72d",
   362 => x"8bb404b5",
   363 => x"b408b5e0",
   364 => x"1381b72d",
   365 => x"8115558b",
   366 => x"7625ffaa",
   367 => x"38029805",
   368 => x"0d0402fc",
   369 => x"050d7251",
   370 => x"70fd2ead",
   371 => x"3870fd24",
   372 => x"8a3870fc",
   373 => x"2e80c438",
   374 => x"8ca30470",
   375 => x"fe2eb138",
   376 => x"70ff2e09",
   377 => x"8106bc38",
   378 => x"b4e40851",
   379 => x"70802eb3",
   380 => x"38ff11b4",
   381 => x"e40c8ca3",
   382 => x"04b4e408",
   383 => x"f00570b4",
   384 => x"e40c5170",
   385 => x"80259c38",
   386 => x"800bb4e4",
   387 => x"0c8ca304",
   388 => x"b4e40881",
   389 => x"05b4e40c",
   390 => x"8ca304b4",
   391 => x"e4089005",
   392 => x"b4e40c8a",
   393 => x"a72da5eb",
   394 => x"2d028405",
   395 => x"0d0402fc",
   396 => x"050d800b",
   397 => x"b4e40c8a",
   398 => x"a72db3b0",
   399 => x"51a7862d",
   400 => x"0284050d",
   401 => x"0402f405",
   402 => x"0d805186",
   403 => x"922d810b",
   404 => x"fec40c80",
   405 => x"0bfec00c",
   406 => x"840bfec4",
   407 => x"0c830bfe",
   408 => x"cc0ca2f6",
   409 => x"2da5892d",
   410 => x"a2db2da2",
   411 => x"db2d81f7",
   412 => x"2d815184",
   413 => x"e52da2db",
   414 => x"2da2db2d",
   415 => x"815184e5",
   416 => x"2db0f051",
   417 => x"85f12d84",
   418 => x"529ced2d",
   419 => x"8ef72db5",
   420 => x"b408802e",
   421 => x"8638fe52",
   422 => x"8da304ff",
   423 => x"12527180",
   424 => x"24e73871",
   425 => x"802e8181",
   426 => x"3886c22d",
   427 => x"b1885187",
   428 => x"e42db5b4",
   429 => x"08802e8f",
   430 => x"38b2c051",
   431 => x"a7862d80",
   432 => x"5184e52d",
   433 => x"8dd104b5",
   434 => x"b408518c",
   435 => x"ae2da595",
   436 => x"2da38e2d",
   437 => x"a7962db5",
   438 => x"b408bc94",
   439 => x"08882bbc",
   440 => x"980807fe",
   441 => x"d80c5386",
   442 => x"ef2db5b4",
   443 => x"08b5d008",
   444 => x"2ea238b5",
   445 => x"b408b5d0",
   446 => x"0cb5b408",
   447 => x"fec00c84",
   448 => x"52725184",
   449 => x"e52da2db",
   450 => x"2da2db2d",
   451 => x"ff125271",
   452 => x"8025ee38",
   453 => x"72802e89",
   454 => x"388a0bfe",
   455 => x"c40c8dd1",
   456 => x"04820bfe",
   457 => x"c40c8dd1",
   458 => x"04b19451",
   459 => x"85f12d80",
   460 => x"0bb5b40c",
   461 => x"028c050d",
   462 => x"0402e805",
   463 => x"0d77797b",
   464 => x"58555580",
   465 => x"53727625",
   466 => x"a3387470",
   467 => x"81055680",
   468 => x"f52d7470",
   469 => x"81055680",
   470 => x"f52d5252",
   471 => x"71712e86",
   472 => x"3881518e",
   473 => x"ee048113",
   474 => x"538ec504",
   475 => x"805170b5",
   476 => x"b40c0298",
   477 => x"050d0402",
   478 => x"d8050d80",
   479 => x"0bbbb80c",
   480 => x"b7b05280",
   481 => x"519fd52d",
   482 => x"b5b40854",
   483 => x"b5b4088c",
   484 => x"38b1a851",
   485 => x"85f12d73",
   486 => x"55949204",
   487 => x"8056810b",
   488 => x"bbdc0c88",
   489 => x"53b1b452",
   490 => x"b7e6518e",
   491 => x"b92db5b4",
   492 => x"08762e09",
   493 => x"81068738",
   494 => x"b5b408bb",
   495 => x"dc0c8853",
   496 => x"b1c052b8",
   497 => x"82518eb9",
   498 => x"2db5b408",
   499 => x"8738b5b4",
   500 => x"08bbdc0c",
   501 => x"bbdc0880",
   502 => x"2e80f638",
   503 => x"baf60b80",
   504 => x"f52dbaf7",
   505 => x"0b80f52d",
   506 => x"71982b71",
   507 => x"902b07ba",
   508 => x"f80b80f5",
   509 => x"2d70882b",
   510 => x"7207baf9",
   511 => x"0b80f52d",
   512 => x"7107bbae",
   513 => x"0b80f52d",
   514 => x"bbaf0b80",
   515 => x"f52d7188",
   516 => x"2b07535f",
   517 => x"54525a56",
   518 => x"57557381",
   519 => x"abaa2e09",
   520 => x"81068d38",
   521 => x"7551a0f5",
   522 => x"2db5b408",
   523 => x"5690bd04",
   524 => x"7382d4d5",
   525 => x"2e8738b1",
   526 => x"cc5190fe",
   527 => x"04b7b052",
   528 => x"75519fd5",
   529 => x"2db5b408",
   530 => x"55b5b408",
   531 => x"802e83c2",
   532 => x"388853b1",
   533 => x"c052b882",
   534 => x"518eb92d",
   535 => x"b5b40889",
   536 => x"38810bbb",
   537 => x"b80c9184",
   538 => x"048853b1",
   539 => x"b452b7e6",
   540 => x"518eb92d",
   541 => x"b5b40880",
   542 => x"2e8a38b1",
   543 => x"e05185f1",
   544 => x"2d91de04",
   545 => x"bbae0b80",
   546 => x"f52d5473",
   547 => x"80d52e09",
   548 => x"810680ca",
   549 => x"38bbaf0b",
   550 => x"80f52d54",
   551 => x"7381aa2e",
   552 => x"098106ba",
   553 => x"38800bb7",
   554 => x"b00b80f5",
   555 => x"2d565474",
   556 => x"81e92e83",
   557 => x"38815474",
   558 => x"81eb2e8c",
   559 => x"38805573",
   560 => x"752e0981",
   561 => x"0682cb38",
   562 => x"b7bb0b80",
   563 => x"f52d5574",
   564 => x"8d38b7bc",
   565 => x"0b80f52d",
   566 => x"5473822e",
   567 => x"86388055",
   568 => x"949204b7",
   569 => x"bd0b80f5",
   570 => x"2d70bbb0",
   571 => x"0cff05bb",
   572 => x"b40cb7be",
   573 => x"0b80f52d",
   574 => x"b7bf0b80",
   575 => x"f52d5876",
   576 => x"05778280",
   577 => x"290570bb",
   578 => x"c00cb7c0",
   579 => x"0b80f52d",
   580 => x"70bbd40c",
   581 => x"bbb80859",
   582 => x"57587680",
   583 => x"2e81a338",
   584 => x"8853b1c0",
   585 => x"52b88251",
   586 => x"8eb92db5",
   587 => x"b40881e2",
   588 => x"38bbb008",
   589 => x"70842bbb",
   590 => x"bc0c70bb",
   591 => x"d00cb7d5",
   592 => x"0b80f52d",
   593 => x"b7d40b80",
   594 => x"f52d7182",
   595 => x"802905b7",
   596 => x"d60b80f5",
   597 => x"2d708480",
   598 => x"802912b7",
   599 => x"d70b80f5",
   600 => x"2d708180",
   601 => x"0a291270",
   602 => x"bbd80cbb",
   603 => x"d4087129",
   604 => x"bbc00805",
   605 => x"70bbc40c",
   606 => x"b7dd0b80",
   607 => x"f52db7dc",
   608 => x"0b80f52d",
   609 => x"71828029",
   610 => x"05b7de0b",
   611 => x"80f52d70",
   612 => x"84808029",
   613 => x"12b7df0b",
   614 => x"80f52d70",
   615 => x"982b81f0",
   616 => x"0a067205",
   617 => x"70bbc80c",
   618 => x"fe117e29",
   619 => x"7705bbcc",
   620 => x"0c525952",
   621 => x"43545e51",
   622 => x"5259525d",
   623 => x"57595794",
   624 => x"9004b7c2",
   625 => x"0b80f52d",
   626 => x"b7c10b80",
   627 => x"f52d7182",
   628 => x"80290570",
   629 => x"bbbc0c70",
   630 => x"a02983ff",
   631 => x"0570892a",
   632 => x"70bbd00c",
   633 => x"b7c70b80",
   634 => x"f52db7c6",
   635 => x"0b80f52d",
   636 => x"71828029",
   637 => x"0570bbd8",
   638 => x"0c7b7129",
   639 => x"1e70bbcc",
   640 => x"0c7dbbc8",
   641 => x"0c7305bb",
   642 => x"c40c555e",
   643 => x"51515555",
   644 => x"815574b5",
   645 => x"b40c02a8",
   646 => x"050d0402",
   647 => x"ec050d76",
   648 => x"70872c71",
   649 => x"80ff0655",
   650 => x"5654bbb8",
   651 => x"088a3873",
   652 => x"882c7481",
   653 => x"ff065455",
   654 => x"b7b052bb",
   655 => x"c0081551",
   656 => x"9fd52db5",
   657 => x"b40854b5",
   658 => x"b408802e",
   659 => x"b338bbb8",
   660 => x"08802e98",
   661 => x"38728429",
   662 => x"b7b00570",
   663 => x"085253a0",
   664 => x"f52db5b4",
   665 => x"08f00a06",
   666 => x"5394fe04",
   667 => x"7210b7b0",
   668 => x"057080e0",
   669 => x"2d5253a1",
   670 => x"a52db5b4",
   671 => x"08537254",
   672 => x"73b5b40c",
   673 => x"0294050d",
   674 => x"0402ec05",
   675 => x"0d767084",
   676 => x"2cbbcc08",
   677 => x"05718f06",
   678 => x"52555372",
   679 => x"8938b7b0",
   680 => x"5273519f",
   681 => x"d52d72a0",
   682 => x"29b7b005",
   683 => x"54807480",
   684 => x"f52d5455",
   685 => x"72752e83",
   686 => x"38815572",
   687 => x"81e52e93",
   688 => x"3874802e",
   689 => x"8e388b14",
   690 => x"80f52d98",
   691 => x"06537280",
   692 => x"2e833880",
   693 => x"5473b5b4",
   694 => x"0c029405",
   695 => x"0d0402cc",
   696 => x"050d7e60",
   697 => x"5e5a800b",
   698 => x"bbc808bb",
   699 => x"cc08595c",
   700 => x"568058bb",
   701 => x"bc08782e",
   702 => x"81ae3877",
   703 => x"8f06a017",
   704 => x"5754738f",
   705 => x"38b7b052",
   706 => x"76518117",
   707 => x"579fd52d",
   708 => x"b7b05680",
   709 => x"7680f52d",
   710 => x"56547474",
   711 => x"2e833881",
   712 => x"547481e5",
   713 => x"2e80f638",
   714 => x"81707506",
   715 => x"555c7380",
   716 => x"2e80ea38",
   717 => x"8b1680f5",
   718 => x"2d980659",
   719 => x"7880de38",
   720 => x"8b537c52",
   721 => x"75518eb9",
   722 => x"2db5b408",
   723 => x"80cf389c",
   724 => x"160851a0",
   725 => x"f52db5b4",
   726 => x"08841b0c",
   727 => x"9a1680e0",
   728 => x"2d51a1a5",
   729 => x"2db5b408",
   730 => x"b5b40888",
   731 => x"1c0cb5b4",
   732 => x"085555bb",
   733 => x"b808802e",
   734 => x"98389416",
   735 => x"80e02d51",
   736 => x"a1a52db5",
   737 => x"b408902b",
   738 => x"83fff00a",
   739 => x"06701651",
   740 => x"5473881b",
   741 => x"0c787a0c",
   742 => x"7b5497de",
   743 => x"04811858",
   744 => x"bbbc0878",
   745 => x"26fed438",
   746 => x"bbb80880",
   747 => x"2eae387a",
   748 => x"51949b2d",
   749 => x"b5b408b5",
   750 => x"b40880ff",
   751 => x"fffff806",
   752 => x"555b7380",
   753 => x"fffffff8",
   754 => x"2e9238b5",
   755 => x"b408fe05",
   756 => x"bbb00829",
   757 => x"bbc40805",
   758 => x"5795f104",
   759 => x"805473b5",
   760 => x"b40c02b4",
   761 => x"050d0402",
   762 => x"f4050d74",
   763 => x"70088105",
   764 => x"710c7008",
   765 => x"bbb40806",
   766 => x"5353718e",
   767 => x"38881308",
   768 => x"51949b2d",
   769 => x"b5b40888",
   770 => x"140c810b",
   771 => x"b5b40c02",
   772 => x"8c050d04",
   773 => x"02f0050d",
   774 => x"75881108",
   775 => x"fe05bbb0",
   776 => x"0829bbc4",
   777 => x"08117208",
   778 => x"bbb40806",
   779 => x"05795553",
   780 => x"54549fd5",
   781 => x"2d029005",
   782 => x"0d0402f0",
   783 => x"050d7588",
   784 => x"1108fe05",
   785 => x"bbb00829",
   786 => x"bbc40811",
   787 => x"7208bbb4",
   788 => x"08060579",
   789 => x"55535454",
   790 => x"9e952d02",
   791 => x"90050d04",
   792 => x"02f4050d",
   793 => x"d45281ff",
   794 => x"720c7108",
   795 => x"5381ff72",
   796 => x"0c72882b",
   797 => x"83fe8006",
   798 => x"72087081",
   799 => x"ff065152",
   800 => x"5381ff72",
   801 => x"0c727107",
   802 => x"882b7208",
   803 => x"7081ff06",
   804 => x"51525381",
   805 => x"ff720c72",
   806 => x"7107882b",
   807 => x"72087081",
   808 => x"ff067207",
   809 => x"b5b40c52",
   810 => x"53028c05",
   811 => x"0d0402f4",
   812 => x"050d7476",
   813 => x"7181ff06",
   814 => x"d40c5353",
   815 => x"bbe00885",
   816 => x"3871892b",
   817 => x"5271982a",
   818 => x"d40c7190",
   819 => x"2a7081ff",
   820 => x"06d40c51",
   821 => x"71882a70",
   822 => x"81ff06d4",
   823 => x"0c517181",
   824 => x"ff06d40c",
   825 => x"72902a70",
   826 => x"81ff06d4",
   827 => x"0c51d408",
   828 => x"7081ff06",
   829 => x"515182b8",
   830 => x"bf527081",
   831 => x"ff2e0981",
   832 => x"06943881",
   833 => x"ff0bd40c",
   834 => x"d4087081",
   835 => x"ff06ff14",
   836 => x"54515171",
   837 => x"e53870b5",
   838 => x"b40c028c",
   839 => x"050d0402",
   840 => x"fc050d81",
   841 => x"c75181ff",
   842 => x"0bd40cff",
   843 => x"11517080",
   844 => x"25f43802",
   845 => x"84050d04",
   846 => x"02f0050d",
   847 => x"9a9f2d8f",
   848 => x"cf538052",
   849 => x"87fc80f7",
   850 => x"5199ae2d",
   851 => x"b5b40854",
   852 => x"b5b40881",
   853 => x"2e098106",
   854 => x"a33881ff",
   855 => x"0bd40c82",
   856 => x"0a52849c",
   857 => x"80e95199",
   858 => x"ae2db5b4",
   859 => x"088b3881",
   860 => x"ff0bd40c",
   861 => x"73539b82",
   862 => x"049a9f2d",
   863 => x"ff135372",
   864 => x"c13872b5",
   865 => x"b40c0290",
   866 => x"050d0402",
   867 => x"f4050d81",
   868 => x"ff0bd40c",
   869 => x"93538052",
   870 => x"87fc80c1",
   871 => x"5199ae2d",
   872 => x"b5b4088b",
   873 => x"3881ff0b",
   874 => x"d40c8153",
   875 => x"9bb8049a",
   876 => x"9f2dff13",
   877 => x"5372df38",
   878 => x"72b5b40c",
   879 => x"028c050d",
   880 => x"0402f005",
   881 => x"0d9a9f2d",
   882 => x"83aa5284",
   883 => x"9c80c851",
   884 => x"99ae2db5",
   885 => x"b408812e",
   886 => x"09810692",
   887 => x"3898e02d",
   888 => x"b5b40883",
   889 => x"ffff0653",
   890 => x"7283aa2e",
   891 => x"97389b8b",
   892 => x"2d9bff04",
   893 => x"81549ce4",
   894 => x"04b1ec51",
   895 => x"85f12d80",
   896 => x"549ce404",
   897 => x"81ff0bd4",
   898 => x"0cb1539a",
   899 => x"b82db5b4",
   900 => x"08802e80",
   901 => x"c0388052",
   902 => x"87fc80fa",
   903 => x"5199ae2d",
   904 => x"b5b408b1",
   905 => x"3881ff0b",
   906 => x"d40cd408",
   907 => x"5381ff0b",
   908 => x"d40c81ff",
   909 => x"0bd40c81",
   910 => x"ff0bd40c",
   911 => x"81ff0bd4",
   912 => x"0c72862a",
   913 => x"708106b5",
   914 => x"b4085651",
   915 => x"5372802e",
   916 => x"93389bf4",
   917 => x"0472822e",
   918 => x"ff9f38ff",
   919 => x"135372ff",
   920 => x"aa387254",
   921 => x"73b5b40c",
   922 => x"0290050d",
   923 => x"0402f005",
   924 => x"0d810bbb",
   925 => x"e00c8454",
   926 => x"d008708f",
   927 => x"2a708106",
   928 => x"51515372",
   929 => x"f33872d0",
   930 => x"0c9a9f2d",
   931 => x"b1fc5185",
   932 => x"f12dd008",
   933 => x"708f2a70",
   934 => x"81065151",
   935 => x"5372f338",
   936 => x"810bd00c",
   937 => x"b1538052",
   938 => x"84d480c0",
   939 => x"5199ae2d",
   940 => x"b5b40881",
   941 => x"2ea13872",
   942 => x"822e0981",
   943 => x"068c38b2",
   944 => x"885185f1",
   945 => x"2d80539e",
   946 => x"8c04ff13",
   947 => x"5372d738",
   948 => x"ff145473",
   949 => x"ffa2389b",
   950 => x"c12db5b4",
   951 => x"08bbe00c",
   952 => x"b5b4088b",
   953 => x"38815287",
   954 => x"fc80d051",
   955 => x"99ae2d81",
   956 => x"ff0bd40c",
   957 => x"d008708f",
   958 => x"2a708106",
   959 => x"51515372",
   960 => x"f33872d0",
   961 => x"0c81ff0b",
   962 => x"d40c8153",
   963 => x"72b5b40c",
   964 => x"0290050d",
   965 => x"0402e805",
   966 => x"0d785681",
   967 => x"ff0bd40c",
   968 => x"d008708f",
   969 => x"2a708106",
   970 => x"51515372",
   971 => x"f3388281",
   972 => x"0bd00c81",
   973 => x"ff0bd40c",
   974 => x"775287fc",
   975 => x"80d85199",
   976 => x"ae2db5b4",
   977 => x"08802e8c",
   978 => x"38b2a051",
   979 => x"85f12d81",
   980 => x"539fcc04",
   981 => x"81ff0bd4",
   982 => x"0c81fe0b",
   983 => x"d40c80ff",
   984 => x"55757084",
   985 => x"05570870",
   986 => x"982ad40c",
   987 => x"70902c70",
   988 => x"81ff06d4",
   989 => x"0c547088",
   990 => x"2c7081ff",
   991 => x"06d40c54",
   992 => x"7081ff06",
   993 => x"d40c54ff",
   994 => x"15557480",
   995 => x"25d33881",
   996 => x"ff0bd40c",
   997 => x"81ff0bd4",
   998 => x"0c81ff0b",
   999 => x"d40c868d",
  1000 => x"a05481ff",
  1001 => x"0bd40cd4",
  1002 => x"0881ff06",
  1003 => x"55748738",
  1004 => x"ff145473",
  1005 => x"ed3881ff",
  1006 => x"0bd40cd0",
  1007 => x"08708f2a",
  1008 => x"70810651",
  1009 => x"515372f3",
  1010 => x"3872d00c",
  1011 => x"72b5b40c",
  1012 => x"0298050d",
  1013 => x"0402e805",
  1014 => x"0d785580",
  1015 => x"5681ff0b",
  1016 => x"d40cd008",
  1017 => x"708f2a70",
  1018 => x"81065151",
  1019 => x"5372f338",
  1020 => x"82810bd0",
  1021 => x"0c81ff0b",
  1022 => x"d40c7752",
  1023 => x"87fc80d1",
  1024 => x"5199ae2d",
  1025 => x"80dbc6df",
  1026 => x"54b5b408",
  1027 => x"802e8a38",
  1028 => x"b0cc5185",
  1029 => x"f12da0ec",
  1030 => x"0481ff0b",
  1031 => x"d40cd408",
  1032 => x"7081ff06",
  1033 => x"51537281",
  1034 => x"fe2e0981",
  1035 => x"069d3880",
  1036 => x"ff5398e0",
  1037 => x"2db5b408",
  1038 => x"75708405",
  1039 => x"570cff13",
  1040 => x"53728025",
  1041 => x"ed388156",
  1042 => x"a0d104ff",
  1043 => x"145473c9",
  1044 => x"3881ff0b",
  1045 => x"d40c81ff",
  1046 => x"0bd40cd0",
  1047 => x"08708f2a",
  1048 => x"70810651",
  1049 => x"515372f3",
  1050 => x"3872d00c",
  1051 => x"75b5b40c",
  1052 => x"0298050d",
  1053 => x"0402f405",
  1054 => x"0d747088",
  1055 => x"2a83fe80",
  1056 => x"06707298",
  1057 => x"2a077288",
  1058 => x"2b87fc80",
  1059 => x"80067398",
  1060 => x"2b81f00a",
  1061 => x"06717307",
  1062 => x"07b5b40c",
  1063 => x"56515351",
  1064 => x"028c050d",
  1065 => x"0402f805",
  1066 => x"0d028e05",
  1067 => x"80f52d74",
  1068 => x"882b0770",
  1069 => x"83ffff06",
  1070 => x"b5b40c51",
  1071 => x"0288050d",
  1072 => x"0402fc05",
  1073 => x"0d725180",
  1074 => x"710c800b",
  1075 => x"84120c02",
  1076 => x"84050d04",
  1077 => x"02f0050d",
  1078 => x"75700884",
  1079 => x"12085353",
  1080 => x"53ff5471",
  1081 => x"712ea838",
  1082 => x"a58f2d84",
  1083 => x"13087084",
  1084 => x"29148811",
  1085 => x"70087081",
  1086 => x"ff068418",
  1087 => x"08811187",
  1088 => x"06841a0c",
  1089 => x"53515551",
  1090 => x"5151a589",
  1091 => x"2d715473",
  1092 => x"b5b40c02",
  1093 => x"90050d04",
  1094 => x"02f8050d",
  1095 => x"a58f2de0",
  1096 => x"08708b2a",
  1097 => x"70810651",
  1098 => x"52527080",
  1099 => x"2e9d38bb",
  1100 => x"e4087084",
  1101 => x"29bbec05",
  1102 => x"7381ff06",
  1103 => x"710c5151",
  1104 => x"bbe40881",
  1105 => x"118706bb",
  1106 => x"e40c5180",
  1107 => x"0bbc8c0c",
  1108 => x"a5822da5",
  1109 => x"892d0288",
  1110 => x"050d0402",
  1111 => x"fc050da5",
  1112 => x"8f2d810b",
  1113 => x"bc8c0ca5",
  1114 => x"892dbc8c",
  1115 => x"085170fa",
  1116 => x"38028405",
  1117 => x"0d0402fc",
  1118 => x"050dbbe4",
  1119 => x"51a1c12d",
  1120 => x"a29851a4",
  1121 => x"fe2da4a8",
  1122 => x"2d028405",
  1123 => x"0d0402f4",
  1124 => x"050da490",
  1125 => x"04b5b408",
  1126 => x"81f02e09",
  1127 => x"81068938",
  1128 => x"810bb5a8",
  1129 => x"0ca49004",
  1130 => x"b5b40881",
  1131 => x"e02e0981",
  1132 => x"06893881",
  1133 => x"0bb5ac0c",
  1134 => x"a49004b5",
  1135 => x"b40852b5",
  1136 => x"ac08802e",
  1137 => x"8838b5b4",
  1138 => x"08818005",
  1139 => x"5271842c",
  1140 => x"728f0653",
  1141 => x"53b5a808",
  1142 => x"802e9938",
  1143 => x"728429b4",
  1144 => x"e8057213",
  1145 => x"81712b70",
  1146 => x"09730806",
  1147 => x"730c5153",
  1148 => x"53a48604",
  1149 => x"728429b4",
  1150 => x"e8057213",
  1151 => x"83712b72",
  1152 => x"0807720c",
  1153 => x"5353800b",
  1154 => x"b5ac0c80",
  1155 => x"0bb5a80c",
  1156 => x"bbe451a1",
  1157 => x"d42db5b4",
  1158 => x"08ff24fe",
  1159 => x"f838800b",
  1160 => x"b5b40c02",
  1161 => x"8c050d04",
  1162 => x"02f8050d",
  1163 => x"b4e8528f",
  1164 => x"51807270",
  1165 => x"8405540c",
  1166 => x"ff115170",
  1167 => x"8025f238",
  1168 => x"0288050d",
  1169 => x"0402f005",
  1170 => x"0d7551a5",
  1171 => x"8f2d7082",
  1172 => x"2cfc06b4",
  1173 => x"e8117210",
  1174 => x"9e067108",
  1175 => x"70722a70",
  1176 => x"83068274",
  1177 => x"2b700974",
  1178 => x"06760c54",
  1179 => x"51565753",
  1180 => x"5153a589",
  1181 => x"2d71b5b4",
  1182 => x"0c029005",
  1183 => x"0d047198",
  1184 => x"0c04ffb0",
  1185 => x"08b5b40c",
  1186 => x"04810bff",
  1187 => x"b00c0480",
  1188 => x"0bffb00c",
  1189 => x"0402fc05",
  1190 => x"0d810bb5",
  1191 => x"b00c8151",
  1192 => x"84e52d02",
  1193 => x"84050d04",
  1194 => x"02fc050d",
  1195 => x"800bb5b0",
  1196 => x"0c805184",
  1197 => x"e52d0284",
  1198 => x"050d0402",
  1199 => x"ec050d76",
  1200 => x"54805287",
  1201 => x"0b881580",
  1202 => x"f52d5653",
  1203 => x"74722483",
  1204 => x"38a05372",
  1205 => x"5182ee2d",
  1206 => x"81128b15",
  1207 => x"80f52d54",
  1208 => x"52727225",
  1209 => x"de380294",
  1210 => x"050d0402",
  1211 => x"f0050dbc",
  1212 => x"9c085481",
  1213 => x"f72d800b",
  1214 => x"bca00c73",
  1215 => x"08802e81",
  1216 => x"8038820b",
  1217 => x"b5c80cbc",
  1218 => x"a0088f06",
  1219 => x"b5c40c73",
  1220 => x"08527183",
  1221 => x"2e963871",
  1222 => x"83268938",
  1223 => x"71812eaf",
  1224 => x"38a6ec04",
  1225 => x"71852e9f",
  1226 => x"38a6ec04",
  1227 => x"881480f5",
  1228 => x"2d841508",
  1229 => x"b2b05354",
  1230 => x"5285f12d",
  1231 => x"71842913",
  1232 => x"70085252",
  1233 => x"a6f00473",
  1234 => x"51a5bb2d",
  1235 => x"a6ec04bc",
  1236 => x"90088815",
  1237 => x"082c7081",
  1238 => x"06515271",
  1239 => x"802e8738",
  1240 => x"b2b451a6",
  1241 => x"e904b2b8",
  1242 => x"5185f12d",
  1243 => x"84140851",
  1244 => x"85f12dbc",
  1245 => x"a0088105",
  1246 => x"bca00c8c",
  1247 => x"1454a5fb",
  1248 => x"04029005",
  1249 => x"0d0471bc",
  1250 => x"9c0ca5eb",
  1251 => x"2dbca008",
  1252 => x"ff05bca4",
  1253 => x"0c0402ec",
  1254 => x"050dbc9c",
  1255 => x"085580f8",
  1256 => x"51a4c52d",
  1257 => x"b5b40881",
  1258 => x"2a708106",
  1259 => x"5152719b",
  1260 => x"388751a4",
  1261 => x"c52db5b4",
  1262 => x"08812a70",
  1263 => x"81065152",
  1264 => x"71802eb1",
  1265 => x"38a7cb04",
  1266 => x"a38e2d87",
  1267 => x"51a4c52d",
  1268 => x"b5b408f4",
  1269 => x"38a7db04",
  1270 => x"a38e2d80",
  1271 => x"f851a4c5",
  1272 => x"2db5b408",
  1273 => x"f338b5b0",
  1274 => x"08813270",
  1275 => x"b5b00c70",
  1276 => x"525284e5",
  1277 => x"2d800bbc",
  1278 => x"940c800b",
  1279 => x"bc980cb5",
  1280 => x"b00882dd",
  1281 => x"3880da51",
  1282 => x"a4c52db5",
  1283 => x"b408802e",
  1284 => x"8a38bc94",
  1285 => x"08818007",
  1286 => x"bc940c80",
  1287 => x"d951a4c5",
  1288 => x"2db5b408",
  1289 => x"802e8a38",
  1290 => x"bc940880",
  1291 => x"c007bc94",
  1292 => x"0c819451",
  1293 => x"a4c52db5",
  1294 => x"b408802e",
  1295 => x"8938bc94",
  1296 => x"089007bc",
  1297 => x"940c8191",
  1298 => x"51a4c52d",
  1299 => x"b5b40880",
  1300 => x"2e8938bc",
  1301 => x"9408a007",
  1302 => x"bc940c81",
  1303 => x"f551a4c5",
  1304 => x"2db5b408",
  1305 => x"802e8938",
  1306 => x"bc940881",
  1307 => x"07bc940c",
  1308 => x"81f251a4",
  1309 => x"c52db5b4",
  1310 => x"08802e89",
  1311 => x"38bc9408",
  1312 => x"8207bc94",
  1313 => x"0c81eb51",
  1314 => x"a4c52db5",
  1315 => x"b408802e",
  1316 => x"8938bc94",
  1317 => x"088407bc",
  1318 => x"940c81f4",
  1319 => x"51a4c52d",
  1320 => x"b5b40880",
  1321 => x"2e8938bc",
  1322 => x"94088807",
  1323 => x"bc940c80",
  1324 => x"d851a4c5",
  1325 => x"2db5b408",
  1326 => x"802e8a38",
  1327 => x"bc980881",
  1328 => x"8007bc98",
  1329 => x"0c9251a4",
  1330 => x"c52db5b4",
  1331 => x"08802e8a",
  1332 => x"38bc9808",
  1333 => x"80c007bc",
  1334 => x"980c9451",
  1335 => x"a4c52db5",
  1336 => x"b408802e",
  1337 => x"8938bc98",
  1338 => x"089007bc",
  1339 => x"980c9151",
  1340 => x"a4c52db5",
  1341 => x"b408802e",
  1342 => x"8938bc98",
  1343 => x"08a007bc",
  1344 => x"980c9d51",
  1345 => x"a4c52db5",
  1346 => x"b408802e",
  1347 => x"8938bc98",
  1348 => x"088107bc",
  1349 => x"980c9b51",
  1350 => x"a4c52db5",
  1351 => x"b408802e",
  1352 => x"8938bc98",
  1353 => x"088207bc",
  1354 => x"980c9c51",
  1355 => x"a4c52db5",
  1356 => x"b408802e",
  1357 => x"8938bc98",
  1358 => x"088407bc",
  1359 => x"980ca351",
  1360 => x"a4c52db5",
  1361 => x"b408802e",
  1362 => x"8938bc98",
  1363 => x"088807bc",
  1364 => x"980c81fd",
  1365 => x"51a4c52d",
  1366 => x"81fa51a4",
  1367 => x"c52daf9c",
  1368 => x"0481f551",
  1369 => x"a4c52db5",
  1370 => x"b408812a",
  1371 => x"70810651",
  1372 => x"5271802e",
  1373 => x"af38bca4",
  1374 => x"08527180",
  1375 => x"2e8938ff",
  1376 => x"12bca40c",
  1377 => x"aba404bc",
  1378 => x"a00810bc",
  1379 => x"a0080570",
  1380 => x"84291651",
  1381 => x"52881208",
  1382 => x"802e8938",
  1383 => x"ff518812",
  1384 => x"0852712d",
  1385 => x"81f251a4",
  1386 => x"c52db5b4",
  1387 => x"08812a70",
  1388 => x"81065152",
  1389 => x"71802eb1",
  1390 => x"38bca008",
  1391 => x"ff11bca4",
  1392 => x"08565353",
  1393 => x"73722589",
  1394 => x"388114bc",
  1395 => x"a40cabe9",
  1396 => x"04721013",
  1397 => x"70842916",
  1398 => x"51528812",
  1399 => x"08802e89",
  1400 => x"38fe5188",
  1401 => x"12085271",
  1402 => x"2d81fd51",
  1403 => x"a4c52db5",
  1404 => x"b408812a",
  1405 => x"70810651",
  1406 => x"5271802e",
  1407 => x"8638800b",
  1408 => x"bca40c81",
  1409 => x"fa51a4c5",
  1410 => x"2db5b408",
  1411 => x"812a7081",
  1412 => x"06515271",
  1413 => x"802e8938",
  1414 => x"bca008ff",
  1415 => x"05bca40c",
  1416 => x"bca40870",
  1417 => x"53547380",
  1418 => x"2e8a388c",
  1419 => x"15ff1555",
  1420 => x"55aca604",
  1421 => x"820bb5c8",
  1422 => x"0c718f06",
  1423 => x"b5c40c81",
  1424 => x"eb51a4c5",
  1425 => x"2db5b408",
  1426 => x"812a7081",
  1427 => x"06515271",
  1428 => x"802ead38",
  1429 => x"7408852e",
  1430 => x"098106a4",
  1431 => x"38881580",
  1432 => x"f52dff05",
  1433 => x"52718816",
  1434 => x"81b72d71",
  1435 => x"982b5271",
  1436 => x"80258838",
  1437 => x"800b8816",
  1438 => x"81b72d74",
  1439 => x"51a5bb2d",
  1440 => x"81f451a4",
  1441 => x"c52db5b4",
  1442 => x"08812a70",
  1443 => x"81065152",
  1444 => x"71802eb3",
  1445 => x"38740885",
  1446 => x"2e098106",
  1447 => x"aa388815",
  1448 => x"80f52d81",
  1449 => x"05527188",
  1450 => x"1681b72d",
  1451 => x"7181ff06",
  1452 => x"8b1680f5",
  1453 => x"2d545272",
  1454 => x"72278738",
  1455 => x"72881681",
  1456 => x"b72d7451",
  1457 => x"a5bb2d80",
  1458 => x"da51a4c5",
  1459 => x"2db5b408",
  1460 => x"812a7081",
  1461 => x"06515271",
  1462 => x"802e80ff",
  1463 => x"38bc9c08",
  1464 => x"bca40855",
  1465 => x"5373802e",
  1466 => x"8a388c13",
  1467 => x"ff155553",
  1468 => x"ade50472",
  1469 => x"08527182",
  1470 => x"2ea63871",
  1471 => x"82268938",
  1472 => x"71812ea9",
  1473 => x"38aedb04",
  1474 => x"71832eb1",
  1475 => x"3871842e",
  1476 => x"09810680",
  1477 => x"c6388813",
  1478 => x"0851a786",
  1479 => x"2daedb04",
  1480 => x"bca40851",
  1481 => x"88130852",
  1482 => x"712daedb",
  1483 => x"04810b88",
  1484 => x"14082bbc",
  1485 => x"900832bc",
  1486 => x"900caed8",
  1487 => x"04881380",
  1488 => x"f52d8105",
  1489 => x"8b1480f5",
  1490 => x"2d535471",
  1491 => x"74248338",
  1492 => x"80547388",
  1493 => x"1481b72d",
  1494 => x"a5eb2d80",
  1495 => x"54800bb5",
  1496 => x"c80c738f",
  1497 => x"06b5c40c",
  1498 => x"a05273bc",
  1499 => x"a4082e09",
  1500 => x"81069838",
  1501 => x"bca008ff",
  1502 => x"05743270",
  1503 => x"09810570",
  1504 => x"72079f2a",
  1505 => x"91713151",
  1506 => x"51535371",
  1507 => x"5182ee2d",
  1508 => x"8114548e",
  1509 => x"7425c638",
  1510 => x"b5b00852",
  1511 => x"71b5b40c",
  1512 => x"0294050d",
  1513 => x"04000000",
  1514 => x"00ffffff",
  1515 => x"ff00ffff",
  1516 => x"ffff00ff",
  1517 => x"ffffff00",
  1518 => x"52657365",
  1519 => x"74000000",
  1520 => x"53617665",
  1521 => x"20736574",
  1522 => x"74696e67",
  1523 => x"73000000",
  1524 => x"5363616e",
  1525 => x"6c696e65",
  1526 => x"73000000",
  1527 => x"4c6f6164",
  1528 => x"20524f4d",
  1529 => x"20100000",
  1530 => x"45786974",
  1531 => x"00000000",
  1532 => x"50432045",
  1533 => x"6e67696e",
  1534 => x"65206d6f",
  1535 => x"64650000",
  1536 => x"54757262",
  1537 => x"6f677261",
  1538 => x"66782031",
  1539 => x"36206d6f",
  1540 => x"64650000",
  1541 => x"56474120",
  1542 => x"2d203331",
  1543 => x"4b487a2c",
  1544 => x"20363048",
  1545 => x"7a000000",
  1546 => x"5456202d",
  1547 => x"20343830",
  1548 => x"692c2036",
  1549 => x"30487a00",
  1550 => x"4261636b",
  1551 => x"00000000",
  1552 => x"46504741",
  1553 => x"50434520",
  1554 => x"43464700",
  1555 => x"52656164",
  1556 => x"20666169",
  1557 => x"6c65640a",
  1558 => x"00000000",
  1559 => x"4661696c",
  1560 => x"65640a00",
  1561 => x"4c6f6164",
  1562 => x"696e6720",
  1563 => x"00000000",
  1564 => x"496e6974",
  1565 => x"69616c69",
  1566 => x"7a696e67",
  1567 => x"20534420",
  1568 => x"63617264",
  1569 => x"0a000000",
  1570 => x"424f4f54",
  1571 => x"20202020",
  1572 => x"50434500",
  1573 => x"43617264",
  1574 => x"20696e69",
  1575 => x"74206661",
  1576 => x"696c6564",
  1577 => x"0a000000",
  1578 => x"4d425220",
  1579 => x"6661696c",
  1580 => x"0a000000",
  1581 => x"46415431",
  1582 => x"36202020",
  1583 => x"00000000",
  1584 => x"46415433",
  1585 => x"32202020",
  1586 => x"00000000",
  1587 => x"4e6f2070",
  1588 => x"61727469",
  1589 => x"74696f6e",
  1590 => x"20736967",
  1591 => x"0a000000",
  1592 => x"42616420",
  1593 => x"70617274",
  1594 => x"0a000000",
  1595 => x"53444843",
  1596 => x"20657272",
  1597 => x"6f72210a",
  1598 => x"00000000",
  1599 => x"53442069",
  1600 => x"6e69742e",
  1601 => x"2e2e0a00",
  1602 => x"53442063",
  1603 => x"61726420",
  1604 => x"72657365",
  1605 => x"74206661",
  1606 => x"696c6564",
  1607 => x"210a0000",
  1608 => x"57726974",
  1609 => x"65206661",
  1610 => x"696c6564",
  1611 => x"0a000000",
  1612 => x"16200000",
  1613 => x"14200000",
  1614 => x"15200000",
  1615 => x"00000002",
  1616 => x"00000002",
  1617 => x"000017b8",
  1618 => x"000004ce",
  1619 => x"00000002",
  1620 => x"000017c0",
  1621 => x"000003a2",
  1622 => x"00000003",
  1623 => x"000019a8",
  1624 => x"00000002",
  1625 => x"00000001",
  1626 => x"000017d0",
  1627 => x"00000001",
  1628 => x"00000003",
  1629 => x"000019a0",
  1630 => x"00000002",
  1631 => x"00000002",
  1632 => x"000017dc",
  1633 => x"0000062e",
  1634 => x"00000002",
  1635 => x"000017e8",
  1636 => x"000012a8",
  1637 => x"00000000",
  1638 => x"00000000",
  1639 => x"00000000",
  1640 => x"000017f0",
  1641 => x"00001800",
  1642 => x"00001814",
  1643 => x"00001828",
  1644 => x"00000002",
  1645 => x"00001ae0",
  1646 => x"000004e3",
  1647 => x"00000002",
  1648 => x"00001af0",
  1649 => x"000004e3",
  1650 => x"00000002",
  1651 => x"00001b00",
  1652 => x"000004e3",
  1653 => x"00000002",
  1654 => x"00001b10",
  1655 => x"000004e3",
  1656 => x"00000002",
  1657 => x"00001b20",
  1658 => x"000004e3",
  1659 => x"00000002",
  1660 => x"00001b30",
  1661 => x"000004e3",
  1662 => x"00000002",
  1663 => x"00001b40",
  1664 => x"000004e3",
  1665 => x"00000002",
  1666 => x"00001b50",
  1667 => x"000004e3",
  1668 => x"00000002",
  1669 => x"00001b60",
  1670 => x"000004e3",
  1671 => x"00000002",
  1672 => x"00001b70",
  1673 => x"000004e3",
  1674 => x"00000002",
  1675 => x"00001b80",
  1676 => x"000004e3",
  1677 => x"00000002",
  1678 => x"00001b90",
  1679 => x"000004e3",
  1680 => x"00000002",
  1681 => x"00001ba0",
  1682 => x"000004e3",
  1683 => x"00000004",
  1684 => x"00001838",
  1685 => x"00001940",
  1686 => x"00000000",
  1687 => x"00000000",
  1688 => x"000005c2",
  1689 => x"00000000",
  1690 => x"00000000",
  1691 => x"00000000",
  1692 => x"00000000",
  1693 => x"00000000",
  1694 => x"00000000",
  1695 => x"00000000",
  1696 => x"00000000",
  1697 => x"00000000",
  1698 => x"00000000",
  1699 => x"00000000",
  1700 => x"00000000",
  1701 => x"00000000",
  1702 => x"00000000",
  1703 => x"00000000",
  1704 => x"00000000",
  1705 => x"00000000",
  1706 => x"00000000",
  1707 => x"00000000",
  1708 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

