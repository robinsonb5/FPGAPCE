-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0baf",
     9 => x"bc080b0b",
    10 => x"0bafc008",
    11 => x"0b0b0baf",
    12 => x"c4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"afc40c0b",
    16 => x"0b0bafc0",
    17 => x"0c0b0b0b",
    18 => x"afbc0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba990",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"afbc70b6",
    57 => x"a8278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"88cf0402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"afcc0c9f",
    65 => x"0bafd00c",
    66 => x"a0717081",
    67 => x"055334af",
    68 => x"d008ff05",
    69 => x"afd00caf",
    70 => x"d0088025",
    71 => x"eb38afcc",
    72 => x"08ff05af",
    73 => x"cc0cafcc",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bafcc",
    94 => x"08258f38",
    95 => x"82b22daf",
    96 => x"cc08ff05",
    97 => x"afcc0c82",
    98 => x"f404afcc",
    99 => x"08afd008",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38afcc08",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134af",
   108 => x"d0088105",
   109 => x"afd00caf",
   110 => x"d008519f",
   111 => x"7125e238",
   112 => x"800bafd0",
   113 => x"0cafcc08",
   114 => x"8105afcc",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"afd00881",
   120 => x"05afd00c",
   121 => x"afd008a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"afd00caf",
   125 => x"cc088105",
   126 => x"afcc0c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800baf",
   155 => x"d40cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bafd4",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"afd40884",
   167 => x"07afd40c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0bac",
   172 => x"c80c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2cafd408",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02f4050d",
   198 => x"74708206",
   199 => x"b6980cac",
   200 => x"e4718106",
   201 => x"54545171",
   202 => x"881481b7",
   203 => x"2d70822a",
   204 => x"70810651",
   205 => x"51709414",
   206 => x"81b72d70",
   207 => x"afbc0c02",
   208 => x"8c050d04",
   209 => x"02f4050d",
   210 => x"aaa852af",
   211 => x"dc519397",
   212 => x"2dafbc08",
   213 => x"802e9538",
   214 => x"b1b852af",
   215 => x"dc5195cd",
   216 => x"2db1b808",
   217 => x"70fec00c",
   218 => x"5186942d",
   219 => x"028c050d",
   220 => x"0402f805",
   221 => x"0db69808",
   222 => x"8206acec",
   223 => x"0b80f52d",
   224 => x"52527080",
   225 => x"2e853871",
   226 => x"810752ac",
   227 => x"f80b80f5",
   228 => x"2d517080",
   229 => x"2e853871",
   230 => x"84075271",
   231 => x"afbc0c02",
   232 => x"88050d04",
   233 => x"02f0050d",
   234 => x"86f12daf",
   235 => x"bc08aaa8",
   236 => x"53afdc52",
   237 => x"5393972d",
   238 => x"afbc0880",
   239 => x"2ea33872",
   240 => x"b1b80cb1",
   241 => x"bc5480fd",
   242 => x"53807470",
   243 => x"8405560c",
   244 => x"ff135372",
   245 => x"8025f238",
   246 => x"b1b852af",
   247 => x"dc5195f3",
   248 => x"2d029005",
   249 => x"0d04a2c9",
   250 => x"2d040402",
   251 => x"e8050d80",
   252 => x"705755b5",
   253 => x"c408752e",
   254 => x"80ca3874",
   255 => x"5192cb2d",
   256 => x"afbc0880",
   257 => x"2eae3875",
   258 => x"9029afe8",
   259 => x"058117af",
   260 => x"bc085657",
   261 => x"528a5373",
   262 => x"70810555",
   263 => x"80f52d72",
   264 => x"70810554",
   265 => x"81b72dff",
   266 => x"13537280",
   267 => x"25e93880",
   268 => x"7281b72d",
   269 => x"81155575",
   270 => x"8b248938",
   271 => x"b5c40875",
   272 => x"26ffb838",
   273 => x"adbc51a4",
   274 => x"a72d0298",
   275 => x"050d0402",
   276 => x"d4050d80",
   277 => x"5186942d",
   278 => x"810bfec4",
   279 => x"0c800bfe",
   280 => x"c00c840b",
   281 => x"fec40c83",
   282 => x"0bfecc0c",
   283 => x"a0aa2da2",
   284 => x"bd2da08f",
   285 => x"2da08f2d",
   286 => x"81f72d81",
   287 => x"5184e52d",
   288 => x"a08f2da0",
   289 => x"8f2d8151",
   290 => x"84e52daa",
   291 => x"b45185f3",
   292 => x"2d9aa62d",
   293 => x"afbc0880",
   294 => x"2e82cf38",
   295 => x"8cb92daf",
   296 => x"bc0853af",
   297 => x"bc088a38",
   298 => x"aacc5185",
   299 => x"f32d8bf2",
   300 => x"0486c42d",
   301 => x"810bfec4",
   302 => x"0c840bfe",
   303 => x"c40caae0",
   304 => x"52afdc51",
   305 => x"93972daf",
   306 => x"bc08802e",
   307 => x"81c138aa",
   308 => x"ec5185f3",
   309 => x"2dafe008",
   310 => x"57807759",
   311 => x"5a767a2e",
   312 => x"8b38811a",
   313 => x"78812a59",
   314 => x"5a77f738",
   315 => x"f71a779f",
   316 => x"ff06545a",
   317 => x"72802e8b",
   318 => x"38fc8017",
   319 => x"afdc5257",
   320 => x"95a02d80",
   321 => x"772580fa",
   322 => x"38795277",
   323 => x"5184802d",
   324 => x"b1b852af",
   325 => x"dc5195cd",
   326 => x"2dafbc08",
   327 => x"802e80c9",
   328 => x"38b1b85b",
   329 => x"80598ad6",
   330 => x"047a7084",
   331 => x"055c0870",
   332 => x"81ff0671",
   333 => x"882c7081",
   334 => x"ff067390",
   335 => x"2c7081ff",
   336 => x"0675982a",
   337 => x"fec80cfe",
   338 => x"c80c58fe",
   339 => x"c80c57fe",
   340 => x"c80c841a",
   341 => x"5a537653",
   342 => x"84807725",
   343 => x"84388480",
   344 => x"53727924",
   345 => x"c4388af2",
   346 => x"04aafc51",
   347 => x"85f32d8b",
   348 => x"8f04afdc",
   349 => x"5195a02d",
   350 => x"fc801781",
   351 => x"1959578a",
   352 => x"8304820b",
   353 => x"fec40c80",
   354 => x"5184e52d",
   355 => x"8b9504ab",
   356 => x"8c5185f3",
   357 => x"2daccc51",
   358 => x"a4a72da0",
   359 => x"c22da4b7",
   360 => x"2dafbc08",
   361 => x"5486f12d",
   362 => x"afbc08fe",
   363 => x"c00c86f1",
   364 => x"2dafbc08",
   365 => x"afd8082e",
   366 => x"9c38afbc",
   367 => x"08afd80c",
   368 => x"84537351",
   369 => x"84e52da0",
   370 => x"8f2da08f",
   371 => x"2dff1353",
   372 => x"728025ee",
   373 => x"3873802e",
   374 => x"89388a0b",
   375 => x"fec40c8b",
   376 => x"9b04820b",
   377 => x"fec40c8b",
   378 => x"9b04aba0",
   379 => x"5185f32d",
   380 => x"805372af",
   381 => x"bc0c02ac",
   382 => x"050d0402",
   383 => x"e8050d77",
   384 => x"797b5855",
   385 => x"55805372",
   386 => x"7625a338",
   387 => x"74708105",
   388 => x"5680f52d",
   389 => x"74708105",
   390 => x"5680f52d",
   391 => x"52527171",
   392 => x"2e863881",
   393 => x"518cb004",
   394 => x"8113538c",
   395 => x"87048051",
   396 => x"70afbc0c",
   397 => x"0298050d",
   398 => x"0402d805",
   399 => x"0d800bb5",
   400 => x"c00cb1b8",
   401 => x"5280519d",
   402 => x"8e2dafbc",
   403 => x"0854afbc",
   404 => x"088c38ab",
   405 => x"b45185f3",
   406 => x"2d735591",
   407 => x"d4048056",
   408 => x"810bb5e4",
   409 => x"0c8853ab",
   410 => x"c052b1ee",
   411 => x"518bfb2d",
   412 => x"afbc0876",
   413 => x"2e098106",
   414 => x"8738afbc",
   415 => x"08b5e40c",
   416 => x"8853abcc",
   417 => x"52b28a51",
   418 => x"8bfb2daf",
   419 => x"bc088738",
   420 => x"afbc08b5",
   421 => x"e40cb5e4",
   422 => x"08802e80",
   423 => x"f638b4fe",
   424 => x"0b80f52d",
   425 => x"b4ff0b80",
   426 => x"f52d7198",
   427 => x"2b71902b",
   428 => x"07b5800b",
   429 => x"80f52d70",
   430 => x"882b7207",
   431 => x"b5810b80",
   432 => x"f52d7107",
   433 => x"b5b60b80",
   434 => x"f52db5b7",
   435 => x"0b80f52d",
   436 => x"71882b07",
   437 => x"535f5452",
   438 => x"5a565755",
   439 => x"7381abaa",
   440 => x"2e098106",
   441 => x"8d387551",
   442 => x"9ea92daf",
   443 => x"bc08568d",
   444 => x"ff047382",
   445 => x"d4d52e87",
   446 => x"38abd851",
   447 => x"8ec004b1",
   448 => x"b8527551",
   449 => x"9d8e2daf",
   450 => x"bc0855af",
   451 => x"bc08802e",
   452 => x"83c23888",
   453 => x"53abcc52",
   454 => x"b28a518b",
   455 => x"fb2dafbc",
   456 => x"08893881",
   457 => x"0bb5c00c",
   458 => x"8ec60488",
   459 => x"53abc052",
   460 => x"b1ee518b",
   461 => x"fb2dafbc",
   462 => x"08802e8a",
   463 => x"38abec51",
   464 => x"85f32d8f",
   465 => x"a004b5b6",
   466 => x"0b80f52d",
   467 => x"547380d5",
   468 => x"2e098106",
   469 => x"80ca38b5",
   470 => x"b70b80f5",
   471 => x"2d547381",
   472 => x"aa2e0981",
   473 => x"06ba3880",
   474 => x"0bb1b80b",
   475 => x"80f52d56",
   476 => x"547481e9",
   477 => x"2e833881",
   478 => x"547481eb",
   479 => x"2e8c3880",
   480 => x"5573752e",
   481 => x"09810682",
   482 => x"cb38b1c3",
   483 => x"0b80f52d",
   484 => x"55748d38",
   485 => x"b1c40b80",
   486 => x"f52d5473",
   487 => x"822e8638",
   488 => x"805591d4",
   489 => x"04b1c50b",
   490 => x"80f52d70",
   491 => x"b5b80cff",
   492 => x"05b5bc0c",
   493 => x"b1c60b80",
   494 => x"f52db1c7",
   495 => x"0b80f52d",
   496 => x"58760577",
   497 => x"82802905",
   498 => x"70b5c80c",
   499 => x"b1c80b80",
   500 => x"f52d70b5",
   501 => x"dc0cb5c0",
   502 => x"08595758",
   503 => x"76802e81",
   504 => x"a3388853",
   505 => x"abcc52b2",
   506 => x"8a518bfb",
   507 => x"2dafbc08",
   508 => x"81e238b5",
   509 => x"b8087084",
   510 => x"2bb5c40c",
   511 => x"70b5d80c",
   512 => x"b1dd0b80",
   513 => x"f52db1dc",
   514 => x"0b80f52d",
   515 => x"71828029",
   516 => x"05b1de0b",
   517 => x"80f52d70",
   518 => x"84808029",
   519 => x"12b1df0b",
   520 => x"80f52d70",
   521 => x"81800a29",
   522 => x"1270b5e0",
   523 => x"0cb5dc08",
   524 => x"7129b5c8",
   525 => x"080570b5",
   526 => x"cc0cb1e5",
   527 => x"0b80f52d",
   528 => x"b1e40b80",
   529 => x"f52d7182",
   530 => x"802905b1",
   531 => x"e60b80f5",
   532 => x"2d708480",
   533 => x"802912b1",
   534 => x"e70b80f5",
   535 => x"2d70982b",
   536 => x"81f00a06",
   537 => x"720570b5",
   538 => x"d00cfe11",
   539 => x"7e297705",
   540 => x"b5d40c52",
   541 => x"59524354",
   542 => x"5e515259",
   543 => x"525d5759",
   544 => x"5791d204",
   545 => x"b1ca0b80",
   546 => x"f52db1c9",
   547 => x"0b80f52d",
   548 => x"71828029",
   549 => x"0570b5c4",
   550 => x"0c70a029",
   551 => x"83ff0570",
   552 => x"892a70b5",
   553 => x"d80cb1cf",
   554 => x"0b80f52d",
   555 => x"b1ce0b80",
   556 => x"f52d7182",
   557 => x"80290570",
   558 => x"b5e00c7b",
   559 => x"71291e70",
   560 => x"b5d40c7d",
   561 => x"b5d00c73",
   562 => x"05b5cc0c",
   563 => x"555e5151",
   564 => x"55558155",
   565 => x"74afbc0c",
   566 => x"02a8050d",
   567 => x"0402ec05",
   568 => x"0d767087",
   569 => x"2c7180ff",
   570 => x"06555654",
   571 => x"b5c0088a",
   572 => x"3873882c",
   573 => x"7481ff06",
   574 => x"5455b1b8",
   575 => x"52b5c808",
   576 => x"15519d8e",
   577 => x"2dafbc08",
   578 => x"54afbc08",
   579 => x"802eb338",
   580 => x"b5c00880",
   581 => x"2e983872",
   582 => x"8429b1b8",
   583 => x"05700852",
   584 => x"539ea92d",
   585 => x"afbc08f0",
   586 => x"0a065392",
   587 => x"c0047210",
   588 => x"b1b80570",
   589 => x"80e02d52",
   590 => x"539ed92d",
   591 => x"afbc0853",
   592 => x"725473af",
   593 => x"bc0c0294",
   594 => x"050d0402",
   595 => x"ec050d76",
   596 => x"70842cb5",
   597 => x"d4080555",
   598 => x"8f065574",
   599 => x"8938b1b8",
   600 => x"5273519d",
   601 => x"8e2d800b",
   602 => x"b1b80b80",
   603 => x"f52d5553",
   604 => x"73732e83",
   605 => x"38815373",
   606 => x"81e52e8e",
   607 => x"3874a029",
   608 => x"b1b80554",
   609 => x"72883893",
   610 => x"8c048053",
   611 => x"725473af",
   612 => x"bc0c0294",
   613 => x"050d0402",
   614 => x"cc050d7e",
   615 => x"605e5a80",
   616 => x"0bb5d008",
   617 => x"b5d40859",
   618 => x"5c568058",
   619 => x"b5c40878",
   620 => x"2e81ae38",
   621 => x"778f06a0",
   622 => x"17575473",
   623 => x"8f38b1b8",
   624 => x"52765181",
   625 => x"17579d8e",
   626 => x"2db1b856",
   627 => x"807680f5",
   628 => x"2d565474",
   629 => x"742e8338",
   630 => x"81547481",
   631 => x"e52e80f6",
   632 => x"38817075",
   633 => x"06555c73",
   634 => x"802e80ea",
   635 => x"388b1680",
   636 => x"f52d9806",
   637 => x"597880de",
   638 => x"388b537c",
   639 => x"5275518b",
   640 => x"fb2dafbc",
   641 => x"0880cf38",
   642 => x"9c160851",
   643 => x"9ea92daf",
   644 => x"bc08841b",
   645 => x"0c9a1680",
   646 => x"e02d519e",
   647 => x"d92dafbc",
   648 => x"08afbc08",
   649 => x"881c0caf",
   650 => x"bc085555",
   651 => x"b5c00880",
   652 => x"2e983894",
   653 => x"1680e02d",
   654 => x"519ed92d",
   655 => x"afbc0890",
   656 => x"2b83fff0",
   657 => x"0a067016",
   658 => x"51547388",
   659 => x"1b0c787a",
   660 => x"0c7b5495",
   661 => x"97048118",
   662 => x"58b5c408",
   663 => x"7826fed4",
   664 => x"38b5c008",
   665 => x"802eae38",
   666 => x"7a5191dd",
   667 => x"2dafbc08",
   668 => x"afbc0880",
   669 => x"fffffff8",
   670 => x"06555b73",
   671 => x"80ffffff",
   672 => x"f82e9238",
   673 => x"afbc08fe",
   674 => x"05b5b808",
   675 => x"29b5cc08",
   676 => x"055793aa",
   677 => x"04805473",
   678 => x"afbc0c02",
   679 => x"b4050d04",
   680 => x"02f4050d",
   681 => x"74700881",
   682 => x"05710c70",
   683 => x"08b5bc08",
   684 => x"06535371",
   685 => x"8e388813",
   686 => x"085191dd",
   687 => x"2dafbc08",
   688 => x"88140c81",
   689 => x"0bafbc0c",
   690 => x"028c050d",
   691 => x"0402f005",
   692 => x"0d758811",
   693 => x"08fe05b5",
   694 => x"b80829b5",
   695 => x"cc081172",
   696 => x"08b5bc08",
   697 => x"06057955",
   698 => x"5354549d",
   699 => x"8e2d0290",
   700 => x"050d0402",
   701 => x"f0050d75",
   702 => x"881108fe",
   703 => x"05b5b808",
   704 => x"29b5cc08",
   705 => x"117208b5",
   706 => x"bc080605",
   707 => x"79555354",
   708 => x"549bce2d",
   709 => x"0290050d",
   710 => x"0402f405",
   711 => x"0dd45281",
   712 => x"ff720c71",
   713 => x"085381ff",
   714 => x"720c7288",
   715 => x"2b83fe80",
   716 => x"06720870",
   717 => x"81ff0651",
   718 => x"525381ff",
   719 => x"720c7271",
   720 => x"07882b72",
   721 => x"087081ff",
   722 => x"06515253",
   723 => x"81ff720c",
   724 => x"72710788",
   725 => x"2b720870",
   726 => x"81ff0672",
   727 => x"07afbc0c",
   728 => x"5253028c",
   729 => x"050d0402",
   730 => x"f4050d74",
   731 => x"767181ff",
   732 => x"06d40c53",
   733 => x"53b5e808",
   734 => x"85387189",
   735 => x"2b527198",
   736 => x"2ad40c71",
   737 => x"902a7081",
   738 => x"ff06d40c",
   739 => x"5171882a",
   740 => x"7081ff06",
   741 => x"d40c5171",
   742 => x"81ff06d4",
   743 => x"0c72902a",
   744 => x"7081ff06",
   745 => x"d40c51d4",
   746 => x"087081ff",
   747 => x"06515182",
   748 => x"b8bf5270",
   749 => x"81ff2e09",
   750 => x"81069438",
   751 => x"81ff0bd4",
   752 => x"0cd40870",
   753 => x"81ff06ff",
   754 => x"14545151",
   755 => x"71e53870",
   756 => x"afbc0c02",
   757 => x"8c050d04",
   758 => x"02fc050d",
   759 => x"81c75181",
   760 => x"ff0bd40c",
   761 => x"ff115170",
   762 => x"8025f438",
   763 => x"0284050d",
   764 => x"0402f005",
   765 => x"0d97d82d",
   766 => x"8fcf5380",
   767 => x"5287fc80",
   768 => x"f75196e7",
   769 => x"2dafbc08",
   770 => x"54afbc08",
   771 => x"812e0981",
   772 => x"06a33881",
   773 => x"ff0bd40c",
   774 => x"820a5284",
   775 => x"9c80e951",
   776 => x"96e72daf",
   777 => x"bc088b38",
   778 => x"81ff0bd4",
   779 => x"0c735398",
   780 => x"bb0497d8",
   781 => x"2dff1353",
   782 => x"72c13872",
   783 => x"afbc0c02",
   784 => x"90050d04",
   785 => x"02f4050d",
   786 => x"81ff0bd4",
   787 => x"0c935380",
   788 => x"5287fc80",
   789 => x"c15196e7",
   790 => x"2dafbc08",
   791 => x"8b3881ff",
   792 => x"0bd40c81",
   793 => x"5398f104",
   794 => x"97d82dff",
   795 => x"135372df",
   796 => x"3872afbc",
   797 => x"0c028c05",
   798 => x"0d0402f0",
   799 => x"050d97d8",
   800 => x"2d83aa52",
   801 => x"849c80c8",
   802 => x"5196e72d",
   803 => x"afbc0881",
   804 => x"2e098106",
   805 => x"92389699",
   806 => x"2dafbc08",
   807 => x"83ffff06",
   808 => x"537283aa",
   809 => x"2e973898",
   810 => x"c42d99b8",
   811 => x"0481549a",
   812 => x"9d04abf8",
   813 => x"5185f32d",
   814 => x"80549a9d",
   815 => x"0481ff0b",
   816 => x"d40cb153",
   817 => x"97f12daf",
   818 => x"bc08802e",
   819 => x"80c03880",
   820 => x"5287fc80",
   821 => x"fa5196e7",
   822 => x"2dafbc08",
   823 => x"b13881ff",
   824 => x"0bd40cd4",
   825 => x"085381ff",
   826 => x"0bd40c81",
   827 => x"ff0bd40c",
   828 => x"81ff0bd4",
   829 => x"0c81ff0b",
   830 => x"d40c7286",
   831 => x"2a708106",
   832 => x"afbc0856",
   833 => x"51537280",
   834 => x"2e933899",
   835 => x"ad047282",
   836 => x"2eff9f38",
   837 => x"ff135372",
   838 => x"ffaa3872",
   839 => x"5473afbc",
   840 => x"0c029005",
   841 => x"0d0402f0",
   842 => x"050d810b",
   843 => x"b5e80c84",
   844 => x"54d00870",
   845 => x"8f2a7081",
   846 => x"06515153",
   847 => x"72f33872",
   848 => x"d00c97d8",
   849 => x"2dac8851",
   850 => x"85f32dd0",
   851 => x"08708f2a",
   852 => x"70810651",
   853 => x"515372f3",
   854 => x"38810bd0",
   855 => x"0cb15380",
   856 => x"5284d480",
   857 => x"c05196e7",
   858 => x"2dafbc08",
   859 => x"812ea138",
   860 => x"72822e09",
   861 => x"81068c38",
   862 => x"ac945185",
   863 => x"f32d8053",
   864 => x"9bc504ff",
   865 => x"135372d7",
   866 => x"38ff1454",
   867 => x"73ffa238",
   868 => x"98fa2daf",
   869 => x"bc08b5e8",
   870 => x"0cafbc08",
   871 => x"8b388152",
   872 => x"87fc80d0",
   873 => x"5196e72d",
   874 => x"81ff0bd4",
   875 => x"0cd00870",
   876 => x"8f2a7081",
   877 => x"06515153",
   878 => x"72f33872",
   879 => x"d00c81ff",
   880 => x"0bd40c81",
   881 => x"5372afbc",
   882 => x"0c029005",
   883 => x"0d0402e8",
   884 => x"050d7856",
   885 => x"81ff0bd4",
   886 => x"0cd00870",
   887 => x"8f2a7081",
   888 => x"06515153",
   889 => x"72f33882",
   890 => x"810bd00c",
   891 => x"81ff0bd4",
   892 => x"0c775287",
   893 => x"fc80d851",
   894 => x"96e72daf",
   895 => x"bc08802e",
   896 => x"8c38acac",
   897 => x"5185f32d",
   898 => x"81539d85",
   899 => x"0481ff0b",
   900 => x"d40c81fe",
   901 => x"0bd40c80",
   902 => x"ff557570",
   903 => x"84055708",
   904 => x"70982ad4",
   905 => x"0c70902c",
   906 => x"7081ff06",
   907 => x"d40c5470",
   908 => x"882c7081",
   909 => x"ff06d40c",
   910 => x"547081ff",
   911 => x"06d40c54",
   912 => x"ff155574",
   913 => x"8025d338",
   914 => x"81ff0bd4",
   915 => x"0c81ff0b",
   916 => x"d40c81ff",
   917 => x"0bd40c86",
   918 => x"8da05481",
   919 => x"ff0bd40c",
   920 => x"d40881ff",
   921 => x"06557487",
   922 => x"38ff1454",
   923 => x"73ed3881",
   924 => x"ff0bd40c",
   925 => x"d008708f",
   926 => x"2a708106",
   927 => x"51515372",
   928 => x"f33872d0",
   929 => x"0c72afbc",
   930 => x"0c029805",
   931 => x"0d0402e8",
   932 => x"050d7855",
   933 => x"805681ff",
   934 => x"0bd40cd0",
   935 => x"08708f2a",
   936 => x"70810651",
   937 => x"515372f3",
   938 => x"3882810b",
   939 => x"d00c81ff",
   940 => x"0bd40c77",
   941 => x"5287fc80",
   942 => x"d15196e7",
   943 => x"2d80dbc6",
   944 => x"df54afbc",
   945 => x"08802e8a",
   946 => x"38aafc51",
   947 => x"85f32d9e",
   948 => x"a00481ff",
   949 => x"0bd40cd4",
   950 => x"087081ff",
   951 => x"06515372",
   952 => x"81fe2e09",
   953 => x"81069d38",
   954 => x"80ff5396",
   955 => x"992dafbc",
   956 => x"08757084",
   957 => x"05570cff",
   958 => x"13537280",
   959 => x"25ed3881",
   960 => x"569e8a04",
   961 => x"ff145473",
   962 => x"c93881ff",
   963 => x"0bd40cd0",
   964 => x"08708f2a",
   965 => x"70810651",
   966 => x"515372f3",
   967 => x"3872d00c",
   968 => x"75afbc0c",
   969 => x"0298050d",
   970 => x"0402f405",
   971 => x"0d747088",
   972 => x"2a83fe80",
   973 => x"06707298",
   974 => x"2a077288",
   975 => x"2b87fc80",
   976 => x"80067398",
   977 => x"2b81f00a",
   978 => x"06717307",
   979 => x"07afbc0c",
   980 => x"56515351",
   981 => x"028c050d",
   982 => x"0402f805",
   983 => x"0d028e05",
   984 => x"80f52d74",
   985 => x"882b0770",
   986 => x"83ffff06",
   987 => x"afbc0c51",
   988 => x"0288050d",
   989 => x"0402fc05",
   990 => x"0d725180",
   991 => x"710c800b",
   992 => x"84120c02",
   993 => x"84050d04",
   994 => x"02f0050d",
   995 => x"75700884",
   996 => x"12085353",
   997 => x"53ff5471",
   998 => x"712ea838",
   999 => x"a2c32d84",
  1000 => x"13087084",
  1001 => x"29148811",
  1002 => x"70087081",
  1003 => x"ff068418",
  1004 => x"08811187",
  1005 => x"06841a0c",
  1006 => x"53515551",
  1007 => x"5151a2bd",
  1008 => x"2d715473",
  1009 => x"afbc0c02",
  1010 => x"90050d04",
  1011 => x"02f8050d",
  1012 => x"a2c32de0",
  1013 => x"08708b2a",
  1014 => x"70810651",
  1015 => x"52527080",
  1016 => x"2e9d38b5",
  1017 => x"ec087084",
  1018 => x"29b5f405",
  1019 => x"7381ff06",
  1020 => x"710c5151",
  1021 => x"b5ec0881",
  1022 => x"118706b5",
  1023 => x"ec0c5180",
  1024 => x"0bb6940c",
  1025 => x"a2b62da2",
  1026 => x"bd2d0288",
  1027 => x"050d0402",
  1028 => x"fc050da2",
  1029 => x"c32d810b",
  1030 => x"b6940ca2",
  1031 => x"bd2db694",
  1032 => x"085170fa",
  1033 => x"38028405",
  1034 => x"0d0402fc",
  1035 => x"050db5ec",
  1036 => x"519ef52d",
  1037 => x"9fcc51a2",
  1038 => x"b22da1dc",
  1039 => x"2d028405",
  1040 => x"0d0402f4",
  1041 => x"050da1c4",
  1042 => x"04afbc08",
  1043 => x"81f02e09",
  1044 => x"81068938",
  1045 => x"810bafb0",
  1046 => x"0ca1c404",
  1047 => x"afbc0881",
  1048 => x"e02e0981",
  1049 => x"06893881",
  1050 => x"0bafb40c",
  1051 => x"a1c404af",
  1052 => x"bc0852af",
  1053 => x"b408802e",
  1054 => x"8838afbc",
  1055 => x"08818005",
  1056 => x"5271842c",
  1057 => x"728f0653",
  1058 => x"53afb008",
  1059 => x"802e9938",
  1060 => x"728429ae",
  1061 => x"f0057213",
  1062 => x"81712b70",
  1063 => x"09730806",
  1064 => x"730c5153",
  1065 => x"53a1ba04",
  1066 => x"728429ae",
  1067 => x"f0057213",
  1068 => x"83712b72",
  1069 => x"0807720c",
  1070 => x"5353800b",
  1071 => x"afb40c80",
  1072 => x"0bafb00c",
  1073 => x"b5ec519f",
  1074 => x"882dafbc",
  1075 => x"08ff24fe",
  1076 => x"f838800b",
  1077 => x"afbc0c02",
  1078 => x"8c050d04",
  1079 => x"02f8050d",
  1080 => x"aef0528f",
  1081 => x"51807270",
  1082 => x"8405540c",
  1083 => x"ff115170",
  1084 => x"8025f238",
  1085 => x"0288050d",
  1086 => x"0402f005",
  1087 => x"0d7551a2",
  1088 => x"c32d7082",
  1089 => x"2cfc06ae",
  1090 => x"f0117210",
  1091 => x"9e067108",
  1092 => x"70722a70",
  1093 => x"83068274",
  1094 => x"2b700974",
  1095 => x"06760c54",
  1096 => x"51565753",
  1097 => x"5153a2bd",
  1098 => x"2d71afbc",
  1099 => x"0c029005",
  1100 => x"0d047198",
  1101 => x"0c04ffb0",
  1102 => x"08afbc0c",
  1103 => x"04810bff",
  1104 => x"b00c0480",
  1105 => x"0bffb00c",
  1106 => x"0402fc05",
  1107 => x"0d800baf",
  1108 => x"b80c8051",
  1109 => x"84e52d02",
  1110 => x"84050d04",
  1111 => x"02ec050d",
  1112 => x"76548052",
  1113 => x"870b8815",
  1114 => x"80f52d56",
  1115 => x"53747224",
  1116 => x"8338a053",
  1117 => x"725182ee",
  1118 => x"2d81128b",
  1119 => x"1580f52d",
  1120 => x"54527272",
  1121 => x"25de3802",
  1122 => x"94050d04",
  1123 => x"02f0050d",
  1124 => x"b69c0854",
  1125 => x"81f72d80",
  1126 => x"0bb6a00c",
  1127 => x"7308802e",
  1128 => x"81803882",
  1129 => x"0bafd00c",
  1130 => x"b6a0088f",
  1131 => x"06afcc0c",
  1132 => x"73085271",
  1133 => x"832e9638",
  1134 => x"71832689",
  1135 => x"3871812e",
  1136 => x"af38a48d",
  1137 => x"0471852e",
  1138 => x"9f38a48d",
  1139 => x"04881480",
  1140 => x"f52d8415",
  1141 => x"08acbc53",
  1142 => x"545285f3",
  1143 => x"2d718429",
  1144 => x"13700852",
  1145 => x"52a49104",
  1146 => x"7351a2dc",
  1147 => x"2da48d04",
  1148 => x"b6980888",
  1149 => x"15082c70",
  1150 => x"81065152",
  1151 => x"71802e87",
  1152 => x"38acc051",
  1153 => x"a48a04ac",
  1154 => x"c45185f3",
  1155 => x"2d841408",
  1156 => x"5185f32d",
  1157 => x"b6a00881",
  1158 => x"05b6a00c",
  1159 => x"8c1454a3",
  1160 => x"9c040290",
  1161 => x"050d0471",
  1162 => x"b69c0ca3",
  1163 => x"8c2db6a0",
  1164 => x"08ff05b6",
  1165 => x"a40c0402",
  1166 => x"ec050db6",
  1167 => x"9c085580",
  1168 => x"f851a1f9",
  1169 => x"2dafbc08",
  1170 => x"812a7081",
  1171 => x"06515271",
  1172 => x"9b388751",
  1173 => x"a1f92daf",
  1174 => x"bc08812a",
  1175 => x"70810651",
  1176 => x"5271802e",
  1177 => x"b138a4ec",
  1178 => x"04a0c22d",
  1179 => x"8751a1f9",
  1180 => x"2dafbc08",
  1181 => x"f438a4fc",
  1182 => x"04a0c22d",
  1183 => x"80f851a1",
  1184 => x"f92dafbc",
  1185 => x"08f338af",
  1186 => x"b8088132",
  1187 => x"70afb80c",
  1188 => x"70525284",
  1189 => x"e52dafb8",
  1190 => x"08a23880",
  1191 => x"da51a1f9",
  1192 => x"2d81f551",
  1193 => x"a1f92d81",
  1194 => x"f251a1f9",
  1195 => x"2d81eb51",
  1196 => x"a1f92d81",
  1197 => x"f451a1f9",
  1198 => x"2da98404",
  1199 => x"81f551a1",
  1200 => x"f92dafbc",
  1201 => x"08812a70",
  1202 => x"81065152",
  1203 => x"71802e8f",
  1204 => x"38b6a408",
  1205 => x"5271802e",
  1206 => x"8638ff12",
  1207 => x"b6a40c81",
  1208 => x"f251a1f9",
  1209 => x"2dafbc08",
  1210 => x"812a7081",
  1211 => x"06515271",
  1212 => x"802e9538",
  1213 => x"b6a008ff",
  1214 => x"05b6a408",
  1215 => x"54527272",
  1216 => x"25863881",
  1217 => x"13b6a40c",
  1218 => x"b6a40870",
  1219 => x"53547380",
  1220 => x"2e8a388c",
  1221 => x"15ff1555",
  1222 => x"55a68e04",
  1223 => x"820bafd0",
  1224 => x"0c718f06",
  1225 => x"afcc0c81",
  1226 => x"eb51a1f9",
  1227 => x"2dafbc08",
  1228 => x"812a7081",
  1229 => x"06515271",
  1230 => x"802ead38",
  1231 => x"7408852e",
  1232 => x"098106a4",
  1233 => x"38881580",
  1234 => x"f52dff05",
  1235 => x"52718816",
  1236 => x"81b72d71",
  1237 => x"982b5271",
  1238 => x"80258838",
  1239 => x"800b8816",
  1240 => x"81b72d74",
  1241 => x"51a2dc2d",
  1242 => x"81f451a1",
  1243 => x"f92dafbc",
  1244 => x"08812a70",
  1245 => x"81065152",
  1246 => x"71802eb3",
  1247 => x"38740885",
  1248 => x"2e098106",
  1249 => x"aa388815",
  1250 => x"80f52d81",
  1251 => x"05527188",
  1252 => x"1681b72d",
  1253 => x"7181ff06",
  1254 => x"8b1680f5",
  1255 => x"2d545272",
  1256 => x"72278738",
  1257 => x"72881681",
  1258 => x"b72d7451",
  1259 => x"a2dc2d80",
  1260 => x"da51a1f9",
  1261 => x"2dafbc08",
  1262 => x"812a7081",
  1263 => x"06515271",
  1264 => x"802e80ff",
  1265 => x"38b69c08",
  1266 => x"b6a40855",
  1267 => x"5373802e",
  1268 => x"8a388c13",
  1269 => x"ff155553",
  1270 => x"a7cd0472",
  1271 => x"08527182",
  1272 => x"2ea63871",
  1273 => x"82268938",
  1274 => x"71812ea9",
  1275 => x"38a8c304",
  1276 => x"71832eb1",
  1277 => x"3871842e",
  1278 => x"09810680",
  1279 => x"c6388813",
  1280 => x"0851a4a7",
  1281 => x"2da8c304",
  1282 => x"b6a40851",
  1283 => x"88130852",
  1284 => x"712da8c3",
  1285 => x"04810b88",
  1286 => x"14082bb6",
  1287 => x"980832b6",
  1288 => x"980ca8c0",
  1289 => x"04881380",
  1290 => x"f52d8105",
  1291 => x"8b1480f5",
  1292 => x"2d535471",
  1293 => x"74248338",
  1294 => x"80547388",
  1295 => x"1481b72d",
  1296 => x"a38c2d80",
  1297 => x"54800baf",
  1298 => x"d00c738f",
  1299 => x"06afcc0c",
  1300 => x"a05273b6",
  1301 => x"a4082e09",
  1302 => x"81069838",
  1303 => x"b6a008ff",
  1304 => x"05743270",
  1305 => x"09810570",
  1306 => x"72079f2a",
  1307 => x"91713151",
  1308 => x"51535371",
  1309 => x"5182ee2d",
  1310 => x"8114548e",
  1311 => x"7425c638",
  1312 => x"afb80852",
  1313 => x"71afbc0c",
  1314 => x"0294050d",
  1315 => x"04000000",
  1316 => x"00ffffff",
  1317 => x"ff00ffff",
  1318 => x"ffff00ff",
  1319 => x"ffffff00",
  1320 => x"52657365",
  1321 => x"74000000",
  1322 => x"53617665",
  1323 => x"20736574",
  1324 => x"74696e67",
  1325 => x"73000000",
  1326 => x"5363616e",
  1327 => x"6c696e65",
  1328 => x"73000000",
  1329 => x"4c6f6164",
  1330 => x"20524f4d",
  1331 => x"20100000",
  1332 => x"45786974",
  1333 => x"00000000",
  1334 => x"50432045",
  1335 => x"6e67696e",
  1336 => x"65206d6f",
  1337 => x"64650000",
  1338 => x"54757262",
  1339 => x"6f677261",
  1340 => x"66782031",
  1341 => x"36206d6f",
  1342 => x"64650000",
  1343 => x"56474120",
  1344 => x"2d203331",
  1345 => x"4b487a2c",
  1346 => x"20363048",
  1347 => x"7a000000",
  1348 => x"5456202d",
  1349 => x"20343830",
  1350 => x"692c2036",
  1351 => x"30487a00",
  1352 => x"4261636b",
  1353 => x"00000000",
  1354 => x"46504741",
  1355 => x"50434520",
  1356 => x"43464700",
  1357 => x"496e6974",
  1358 => x"69616c69",
  1359 => x"7a696e67",
  1360 => x"20534420",
  1361 => x"63617264",
  1362 => x"0a000000",
  1363 => x"46696c65",
  1364 => x"73797374",
  1365 => x"656d2065",
  1366 => x"72726f72",
  1367 => x"0a000000",
  1368 => x"4d535833",
  1369 => x"42494f53",
  1370 => x"53595300",
  1371 => x"4c6f6164",
  1372 => x"696e6720",
  1373 => x"524f4d0a",
  1374 => x"00000000",
  1375 => x"52656164",
  1376 => x"20666169",
  1377 => x"6c65640a",
  1378 => x"00000000",
  1379 => x"524f4d20",
  1380 => x"6c6f6164",
  1381 => x"696e6720",
  1382 => x"6661696c",
  1383 => x"65640a00",
  1384 => x"43617264",
  1385 => x"20696e69",
  1386 => x"74206661",
  1387 => x"696c6564",
  1388 => x"0a000000",
  1389 => x"4d425220",
  1390 => x"6661696c",
  1391 => x"0a000000",
  1392 => x"46415431",
  1393 => x"36202020",
  1394 => x"00000000",
  1395 => x"46415433",
  1396 => x"32202020",
  1397 => x"00000000",
  1398 => x"4e6f2070",
  1399 => x"61727469",
  1400 => x"74696f6e",
  1401 => x"20736967",
  1402 => x"0a000000",
  1403 => x"42616420",
  1404 => x"70617274",
  1405 => x"0a000000",
  1406 => x"53444843",
  1407 => x"20657272",
  1408 => x"6f72210a",
  1409 => x"00000000",
  1410 => x"53442069",
  1411 => x"6e69742e",
  1412 => x"2e2e0a00",
  1413 => x"53442063",
  1414 => x"61726420",
  1415 => x"72657365",
  1416 => x"74206661",
  1417 => x"696c6564",
  1418 => x"210a0000",
  1419 => x"57726974",
  1420 => x"65206661",
  1421 => x"696c6564",
  1422 => x"0a000000",
  1423 => x"16200000",
  1424 => x"14200000",
  1425 => x"15200000",
  1426 => x"00000002",
  1427 => x"00000002",
  1428 => x"000014a0",
  1429 => x"000003e6",
  1430 => x"00000002",
  1431 => x"000014a8",
  1432 => x"000003a4",
  1433 => x"00000003",
  1434 => x"000016b4",
  1435 => x"00000002",
  1436 => x"00000001",
  1437 => x"000014b8",
  1438 => x"00000001",
  1439 => x"00000003",
  1440 => x"000016ac",
  1441 => x"00000002",
  1442 => x"00000002",
  1443 => x"000014c4",
  1444 => x"000003eb",
  1445 => x"00000002",
  1446 => x"000014d0",
  1447 => x"00001149",
  1448 => x"00000000",
  1449 => x"00000000",
  1450 => x"00000000",
  1451 => x"000014d8",
  1452 => x"000014e8",
  1453 => x"000014fc",
  1454 => x"00001510",
  1455 => x"00000002",
  1456 => x"000017e8",
  1457 => x"000003ea",
  1458 => x"00000002",
  1459 => x"000017f8",
  1460 => x"000003ea",
  1461 => x"00000002",
  1462 => x"00001808",
  1463 => x"000003ea",
  1464 => x"00000002",
  1465 => x"00001818",
  1466 => x"000003ea",
  1467 => x"00000002",
  1468 => x"00001828",
  1469 => x"000003ea",
  1470 => x"00000002",
  1471 => x"00001838",
  1472 => x"000003ea",
  1473 => x"00000002",
  1474 => x"00001848",
  1475 => x"000003ea",
  1476 => x"00000002",
  1477 => x"00001858",
  1478 => x"000003ea",
  1479 => x"00000002",
  1480 => x"00001868",
  1481 => x"000003ea",
  1482 => x"00000002",
  1483 => x"00001878",
  1484 => x"000003ea",
  1485 => x"00000002",
  1486 => x"00001888",
  1487 => x"000003ea",
  1488 => x"00000002",
  1489 => x"00001898",
  1490 => x"000003ea",
  1491 => x"00000002",
  1492 => x"000018a8",
  1493 => x"000003ea",
  1494 => x"00000004",
  1495 => x"00001520",
  1496 => x"0000164c",
  1497 => x"00000000",
  1498 => x"00000000",
  1499 => x"00000000",
  1500 => x"00000000",
  1501 => x"00000000",
  1502 => x"00000000",
  1503 => x"00000000",
  1504 => x"00000000",
  1505 => x"00000000",
  1506 => x"00000000",
  1507 => x"00000000",
  1508 => x"00000000",
  1509 => x"00000000",
  1510 => x"00000000",
  1511 => x"00000000",
  1512 => x"00000000",
  1513 => x"00000000",
  1514 => x"00000000",
  1515 => x"00000000",
  1516 => x"00000000",
  1517 => x"00000000",
  1518 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

