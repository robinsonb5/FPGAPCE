-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM1 is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM1;

architecture arch of CtrlROM_ROM1 is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b80c2",
     9 => x"b8080b0b",
    10 => x"80c2bc08",
    11 => x"0b0b80c2",
    12 => x"c0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"c2c00c0b",
    16 => x"0b80c2bc",
    17 => x"0c0b0b80",
    18 => x"c2b80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bbc90",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80c2b870",
    57 => x"80ccf827",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c5190c4",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80c2",
    65 => x"c80c9f0b",
    66 => x"80c2cc0c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"c2cc08ff",
    70 => x"0580c2cc",
    71 => x"0c80c2cc",
    72 => x"088025e8",
    73 => x"3880c2c8",
    74 => x"08ff0580",
    75 => x"c2c80c80",
    76 => x"c2c80880",
    77 => x"25d03802",
    78 => x"84050d04",
    79 => x"02f0050d",
    80 => x"f88053f8",
    81 => x"a05483bf",
    82 => x"52737081",
    83 => x"05553351",
    84 => x"70737081",
    85 => x"055534ff",
    86 => x"12527180",
    87 => x"25eb38fb",
    88 => x"c0539f52",
    89 => x"a0737081",
    90 => x"055534ff",
    91 => x"12527180",
    92 => x"25f23802",
    93 => x"90050d04",
    94 => x"02f4050d",
    95 => x"74538e0b",
    96 => x"80c2c808",
    97 => x"25913882",
    98 => x"bc2d80c2",
    99 => x"c808ff05",
   100 => x"80c2c80c",
   101 => x"82fe0480",
   102 => x"c2c80880",
   103 => x"c2cc0853",
   104 => x"51728a2e",
   105 => x"098106be",
   106 => x"38715171",
   107 => x"9f24a438",
   108 => x"80c2c808",
   109 => x"a02911f8",
   110 => x"80115151",
   111 => x"a0713480",
   112 => x"c2cc0881",
   113 => x"0580c2cc",
   114 => x"0c80c2cc",
   115 => x"08519f71",
   116 => x"25de3880",
   117 => x"0b80c2cc",
   118 => x"0c80c2c8",
   119 => x"08810580",
   120 => x"c2c80c83",
   121 => x"fc0470a0",
   122 => x"2912f880",
   123 => x"11515172",
   124 => x"713480c2",
   125 => x"cc088105",
   126 => x"80c2cc0c",
   127 => x"80c2cc08",
   128 => x"a02e0981",
   129 => x"06913880",
   130 => x"0b80c2cc",
   131 => x"0c80c2c8",
   132 => x"08810580",
   133 => x"c2c80c02",
   134 => x"8c050d04",
   135 => x"02e8050d",
   136 => x"77795656",
   137 => x"880bfc16",
   138 => x"77712c8f",
   139 => x"06545254",
   140 => x"80537272",
   141 => x"25953871",
   142 => x"53fbe014",
   143 => x"51877134",
   144 => x"8114ff14",
   145 => x"545472f1",
   146 => x"387153f9",
   147 => x"1576712c",
   148 => x"87065351",
   149 => x"71802e8b",
   150 => x"38fbe014",
   151 => x"51717134",
   152 => x"81145472",
   153 => x"8e249538",
   154 => x"8f733153",
   155 => x"fbe01451",
   156 => x"a0713481",
   157 => x"14ff1454",
   158 => x"5472f138",
   159 => x"0298050d",
   160 => x"0402ec05",
   161 => x"0d800b80",
   162 => x"c2d00cf6",
   163 => x"8c08f690",
   164 => x"0871882c",
   165 => x"565481ff",
   166 => x"06527372",
   167 => x"25893871",
   168 => x"54820b80",
   169 => x"c2d00c72",
   170 => x"882c7381",
   171 => x"ff065455",
   172 => x"7473258d",
   173 => x"387280c2",
   174 => x"d0088407",
   175 => x"80c2d00c",
   176 => x"5573842b",
   177 => x"87e87125",
   178 => x"83713170",
   179 => x"0b0b0bbf",
   180 => x"980c8171",
   181 => x"2bf6880c",
   182 => x"fde813ff",
   183 => x"122c7888",
   184 => x"29ff9405",
   185 => x"70812c80",
   186 => x"c2d00852",
   187 => x"58525551",
   188 => x"52547680",
   189 => x"2e853870",
   190 => x"81075170",
   191 => x"f6940c71",
   192 => x"098105f6",
   193 => x"800c7209",
   194 => x"8105f684",
   195 => x"0c029405",
   196 => x"0d0402f4",
   197 => x"050d7453",
   198 => x"72708105",
   199 => x"5480f52d",
   200 => x"5271802e",
   201 => x"89387151",
   202 => x"82f82d86",
   203 => x"9804028c",
   204 => x"050d0402",
   205 => x"f4050d74",
   206 => x"70820680",
   207 => x"ccdc0cbf",
   208 => x"b4718106",
   209 => x"54545171",
   210 => x"881481b7",
   211 => x"2d70822a",
   212 => x"70810651",
   213 => x"5170a014",
   214 => x"81b72d70",
   215 => x"80c2b80c",
   216 => x"028c050d",
   217 => x"0402f805",
   218 => x"0dbdb052",
   219 => x"80c2d451",
   220 => x"9dd52d80",
   221 => x"c2b80880",
   222 => x"2ea33880",
   223 => x"c5f05280",
   224 => x"c2d451a0",
   225 => x"a22d80c5",
   226 => x"f00880c2",
   227 => x"e00c80c5",
   228 => x"f008fec0",
   229 => x"0c80c5f0",
   230 => x"085186b3",
   231 => x"2d028805",
   232 => x"0d0402f0",
   233 => x"050d8051",
   234 => x"93892dbd",
   235 => x"b05280c2",
   236 => x"d4519dd5",
   237 => x"2d80c2b8",
   238 => x"08802eaa",
   239 => x"3880c2e0",
   240 => x"0880c5f0",
   241 => x"0c80c5f4",
   242 => x"5480fd53",
   243 => x"80747084",
   244 => x"05560cff",
   245 => x"13537280",
   246 => x"25f23880",
   247 => x"c5f05280",
   248 => x"c2d451a0",
   249 => x"cb2d0290",
   250 => x"050d0402",
   251 => x"d4050d80",
   252 => x"c2e008fe",
   253 => x"c00c810b",
   254 => x"fec40c84",
   255 => x"0bfec40c",
   256 => x"7c5280c2",
   257 => x"d4519dd5",
   258 => x"2d80c2b8",
   259 => x"085380c2",
   260 => x"b808802e",
   261 => x"81d43880",
   262 => x"c2d80856",
   263 => x"800bff17",
   264 => x"58597679",
   265 => x"2e8b3881",
   266 => x"1977812a",
   267 => x"585976f7",
   268 => x"38f71976",
   269 => x"9fff0654",
   270 => x"5972802e",
   271 => x"8c38fc80",
   272 => x"1680c2d4",
   273 => x"52569ff2",
   274 => x"2d75b080",
   275 => x"802e0981",
   276 => x"06893882",
   277 => x"0bfedc0c",
   278 => x"88f20475",
   279 => x"9880802e",
   280 => x"09810689",
   281 => x"38810bfe",
   282 => x"dc0c88f2",
   283 => x"04800bfe",
   284 => x"dc0c815b",
   285 => x"80762580",
   286 => x"ef387852",
   287 => x"7651849c",
   288 => x"2d80c5f0",
   289 => x"5280c2d4",
   290 => x"51a0a22d",
   291 => x"80c2b808",
   292 => x"802ebc38",
   293 => x"80c5f05a",
   294 => x"83fc5879",
   295 => x"7084055b",
   296 => x"087083fe",
   297 => x"80067188",
   298 => x"2b83fe80",
   299 => x"0671882a",
   300 => x"0772882a",
   301 => x"83fe8006",
   302 => x"73982a07",
   303 => x"fec80cfe",
   304 => x"c80c56fc",
   305 => x"19595377",
   306 => x"8025d038",
   307 => x"89d70480",
   308 => x"c2b8085b",
   309 => x"84805680",
   310 => x"c2d4519f",
   311 => x"f22dfc80",
   312 => x"16811858",
   313 => x"5688f404",
   314 => x"7a537280",
   315 => x"c2b80c02",
   316 => x"ac050d04",
   317 => x"02fc050d",
   318 => x"adf62dfe",
   319 => x"c4518171",
   320 => x"0c82710c",
   321 => x"0284050d",
   322 => x"0402f405",
   323 => x"0d747678",
   324 => x"53545280",
   325 => x"71259738",
   326 => x"72708105",
   327 => x"5480f52d",
   328 => x"72708105",
   329 => x"5481b72d",
   330 => x"ff115170",
   331 => x"eb388072",
   332 => x"81b72d02",
   333 => x"8c050d04",
   334 => x"02e8050d",
   335 => x"77568070",
   336 => x"56547376",
   337 => x"24b63880",
   338 => x"cc800874",
   339 => x"2eae3873",
   340 => x"519b9a2d",
   341 => x"80c2b808",
   342 => x"80c2b808",
   343 => x"09810570",
   344 => x"80c2b808",
   345 => x"079f2a77",
   346 => x"05811757",
   347 => x"57535374",
   348 => x"76248938",
   349 => x"80cc8008",
   350 => x"7426d438",
   351 => x"7280c2b8",
   352 => x"0c029805",
   353 => x"0d0402f4",
   354 => x"050d80c1",
   355 => x"e4081551",
   356 => x"8ab82d80",
   357 => x"c2b80880",
   358 => x"2e96388b",
   359 => x"5380c2b8",
   360 => x"085280c9",
   361 => x"f0518a89",
   362 => x"2d80c9f0",
   363 => x"5187eb2d",
   364 => x"bf9c51af",
   365 => x"dd2dadf6",
   366 => x"2d805185",
   367 => x"812d028c",
   368 => x"050d0402",
   369 => x"dc050d80",
   370 => x"705a5574",
   371 => x"80c1e408",
   372 => x"25b43880",
   373 => x"cc800875",
   374 => x"2eac3878",
   375 => x"519b9a2d",
   376 => x"80c2b808",
   377 => x"09810570",
   378 => x"80c2b808",
   379 => x"079f2a76",
   380 => x"05811b5b",
   381 => x"56547480",
   382 => x"c1e40825",
   383 => x"893880cc",
   384 => x"80087926",
   385 => x"d6388055",
   386 => x"7880cc80",
   387 => x"082781db",
   388 => x"3878519b",
   389 => x"9a2d80c2",
   390 => x"b808802e",
   391 => x"81ad3880",
   392 => x"c2b8088b",
   393 => x"0580f52d",
   394 => x"70842a70",
   395 => x"81067710",
   396 => x"78842b80",
   397 => x"c9f00b80",
   398 => x"f52d5c5c",
   399 => x"53515556",
   400 => x"73802e80",
   401 => x"cb387416",
   402 => x"822b8e8f",
   403 => x"0b80c0b8",
   404 => x"120c5477",
   405 => x"75311080",
   406 => x"c2e81155",
   407 => x"56907470",
   408 => x"81055681",
   409 => x"b72da074",
   410 => x"81b72d76",
   411 => x"81ff0681",
   412 => x"16585473",
   413 => x"802e8a38",
   414 => x"9c5380c9",
   415 => x"f0528d88",
   416 => x"048b5380",
   417 => x"c2b80852",
   418 => x"80c2ea16",
   419 => x"518dc304",
   420 => x"7416822b",
   421 => x"8b860b80",
   422 => x"c0b8120c",
   423 => x"547681ff",
   424 => x"06811658",
   425 => x"5473802e",
   426 => x"8a389c53",
   427 => x"80c9f052",
   428 => x"8dba048b",
   429 => x"5380c2b8",
   430 => x"08527775",
   431 => x"311080c2",
   432 => x"e8055176",
   433 => x"558a892d",
   434 => x"8de00474",
   435 => x"90297531",
   436 => x"701080c2",
   437 => x"e8055154",
   438 => x"80c2b808",
   439 => x"7481b72d",
   440 => x"81195974",
   441 => x"8b24a338",
   442 => x"8c880474",
   443 => x"90297531",
   444 => x"701080c2",
   445 => x"e8058c77",
   446 => x"31575154",
   447 => x"807481b7",
   448 => x"2d9e14ff",
   449 => x"16565474",
   450 => x"f33802a4",
   451 => x"050d0402",
   452 => x"fc050d80",
   453 => x"c1e40813",
   454 => x"518ab82d",
   455 => x"80c2b808",
   456 => x"802e8938",
   457 => x"80c2b808",
   458 => x"5193892d",
   459 => x"800b80c1",
   460 => x"e40c8bc3",
   461 => x"2daeba2d",
   462 => x"0284050d",
   463 => x"0402fc05",
   464 => x"0d725170",
   465 => x"fd2eb038",
   466 => x"70fd248a",
   467 => x"3870fc2e",
   468 => x"80cc388f",
   469 => x"a80470fe",
   470 => x"2eb73870",
   471 => x"ff2e0981",
   472 => x"0680c538",
   473 => x"80c1e408",
   474 => x"5170802e",
   475 => x"bb38ff11",
   476 => x"80c1e40c",
   477 => x"8fa80480",
   478 => x"c1e408f0",
   479 => x"057080c1",
   480 => x"e40c5170",
   481 => x"8025a138",
   482 => x"800b80c1",
   483 => x"e40c8fa8",
   484 => x"0480c1e4",
   485 => x"08810580",
   486 => x"c1e40c8f",
   487 => x"a80480c1",
   488 => x"e4089005",
   489 => x"80c1e40c",
   490 => x"8bc32dae",
   491 => x"ba2d0284",
   492 => x"050d0402",
   493 => x"fc050d80",
   494 => x"c2e008fb",
   495 => x"0680c2e0",
   496 => x"0c72518b",
   497 => x"862d0284",
   498 => x"050d0402",
   499 => x"fc050d80",
   500 => x"c2e00884",
   501 => x"0780c2e0",
   502 => x"0c72518b",
   503 => x"862d0284",
   504 => x"050d0402",
   505 => x"fc050d80",
   506 => x"0b80c1e4",
   507 => x"0c8bc32d",
   508 => x"80c0b051",
   509 => x"afdd2d80",
   510 => x"c09851af",
   511 => x"f02d0284",
   512 => x"050d0402",
   513 => x"f8050d80",
   514 => x"ccdc0882",
   515 => x"06bfbc0b",
   516 => x"80f52d52",
   517 => x"5270802e",
   518 => x"85387181",
   519 => x"0752bfd4",
   520 => x"0b80f52d",
   521 => x"5170802e",
   522 => x"85387184",
   523 => x"075280c2",
   524 => x"e408802e",
   525 => x"85387190",
   526 => x"07527180",
   527 => x"c2b80c02",
   528 => x"88050d04",
   529 => x"02f4050d",
   530 => x"810b80c2",
   531 => x"e40c9051",
   532 => x"86b32d81",
   533 => x"0bfec40c",
   534 => x"900bfec0",
   535 => x"0c840bfe",
   536 => x"c40c830b",
   537 => x"fecc0cab",
   538 => x"af2dadd6",
   539 => x"2dab922d",
   540 => x"ab922d81",
   541 => x"f92d8151",
   542 => x"85812dab",
   543 => x"922dab92",
   544 => x"2d815185",
   545 => x"812dbdbc",
   546 => x"5186922d",
   547 => x"8452a591",
   548 => x"2d94af2d",
   549 => x"80c2b808",
   550 => x"802e8638",
   551 => x"fe5291a9",
   552 => x"04ff1252",
   553 => x"718024e6",
   554 => x"3871802e",
   555 => x"818b3886",
   556 => x"e52dbdd4",
   557 => x"5187eb2d",
   558 => x"80c2b808",
   559 => x"802e8f38",
   560 => x"bf9c51af",
   561 => x"dd2d8051",
   562 => x"85812d91",
   563 => x"d90480c2",
   564 => x"b808518f",
   565 => x"e32dade2",
   566 => x"2dabc82d",
   567 => x"aff62d80",
   568 => x"c2b80880",
   569 => x"cce00888",
   570 => x"2b80cce4",
   571 => x"0807fed8",
   572 => x"0c539083",
   573 => x"2d80c2b8",
   574 => x"0880c2e0",
   575 => x"082ea538",
   576 => x"80c2b808",
   577 => x"80c2e00c",
   578 => x"80c2b808",
   579 => x"fec00c84",
   580 => x"52725185",
   581 => x"812dab92",
   582 => x"2dab922d",
   583 => x"ff125271",
   584 => x"8025ee38",
   585 => x"72802e89",
   586 => x"388a0bfe",
   587 => x"c40c91d9",
   588 => x"04820bfe",
   589 => x"c40c91d9",
   590 => x"04bde051",
   591 => x"86922d80",
   592 => x"0b80c2b8",
   593 => x"0c028c05",
   594 => x"0d0402e8",
   595 => x"050d7779",
   596 => x"7b585555",
   597 => x"80537276",
   598 => x"25a33874",
   599 => x"70810556",
   600 => x"80f52d74",
   601 => x"70810556",
   602 => x"80f52d52",
   603 => x"5271712e",
   604 => x"86388151",
   605 => x"92ff0481",
   606 => x"135392d6",
   607 => x"04805170",
   608 => x"80c2b80c",
   609 => x"0298050d",
   610 => x"0402ec05",
   611 => x"0d765574",
   612 => x"802e80c2",
   613 => x"389a1580",
   614 => x"e02d51a9",
   615 => x"d52d80c2",
   616 => x"b80880c2",
   617 => x"b80880cc",
   618 => x"a00c80c2",
   619 => x"b8085454",
   620 => x"80cbfc08",
   621 => x"802e9a38",
   622 => x"941580e0",
   623 => x"2d51a9d5",
   624 => x"2d80c2b8",
   625 => x"08902b83",
   626 => x"fff00a06",
   627 => x"70750751",
   628 => x"537280cc",
   629 => x"a00c80cc",
   630 => x"a0085372",
   631 => x"802e9d38",
   632 => x"80cbf408",
   633 => x"fe147129",
   634 => x"80cc8808",
   635 => x"0580cca4",
   636 => x"0c70842b",
   637 => x"80cc800c",
   638 => x"5494aa04",
   639 => x"80cc8c08",
   640 => x"80cca00c",
   641 => x"80cc9008",
   642 => x"80cca40c",
   643 => x"80cbfc08",
   644 => x"802e8b38",
   645 => x"80cbf408",
   646 => x"842b5394",
   647 => x"a50480cc",
   648 => x"9408842b",
   649 => x"537280cc",
   650 => x"800c0294",
   651 => x"050d0402",
   652 => x"d8050d80",
   653 => x"0b80cbfc",
   654 => x"0c80c5f0",
   655 => x"528051a8",
   656 => x"812d80c2",
   657 => x"b8085480",
   658 => x"c2b8088c",
   659 => x"38bdf451",
   660 => x"86922d73",
   661 => x"559a9704",
   662 => x"8056810b",
   663 => x"80cca80c",
   664 => x"8853be80",
   665 => x"5280c6a6",
   666 => x"5192ca2d",
   667 => x"80c2b808",
   668 => x"762e0981",
   669 => x"06893880",
   670 => x"c2b80880",
   671 => x"cca80c88",
   672 => x"53be8c52",
   673 => x"80c6c251",
   674 => x"92ca2d80",
   675 => x"c2b80889",
   676 => x"3880c2b8",
   677 => x"0880cca8",
   678 => x"0c80cca8",
   679 => x"08802e81",
   680 => x"803880c9",
   681 => x"b60b80f5",
   682 => x"2d80c9b7",
   683 => x"0b80f52d",
   684 => x"71982b71",
   685 => x"902b0780",
   686 => x"c9b80b80",
   687 => x"f52d7088",
   688 => x"2b720780",
   689 => x"c9b90b80",
   690 => x"f52d7107",
   691 => x"80c9ee0b",
   692 => x"80f52d80",
   693 => x"c9ef0b80",
   694 => x"f52d7188",
   695 => x"2b07535f",
   696 => x"54525a56",
   697 => x"57557381",
   698 => x"abaa2e09",
   699 => x"81068e38",
   700 => x"7551a9a4",
   701 => x"2d80c2b8",
   702 => x"0856968a",
   703 => x"047382d4",
   704 => x"d52e8738",
   705 => x"be985196",
   706 => x"d30480c5",
   707 => x"f0527551",
   708 => x"a8812d80",
   709 => x"c2b80855",
   710 => x"80c2b808",
   711 => x"802e83f7",
   712 => x"388853be",
   713 => x"8c5280c6",
   714 => x"c25192ca",
   715 => x"2d80c2b8",
   716 => x"088a3881",
   717 => x"0b80cbfc",
   718 => x"0c96d904",
   719 => x"8853be80",
   720 => x"5280c6a6",
   721 => x"5192ca2d",
   722 => x"80c2b808",
   723 => x"802e8a38",
   724 => x"beac5186",
   725 => x"922d97b8",
   726 => x"0480c9ee",
   727 => x"0b80f52d",
   728 => x"547380d5",
   729 => x"2e098106",
   730 => x"80ce3880",
   731 => x"c9ef0b80",
   732 => x"f52d5473",
   733 => x"81aa2e09",
   734 => x"8106bd38",
   735 => x"800b80c5",
   736 => x"f00b80f5",
   737 => x"2d565474",
   738 => x"81e92e83",
   739 => x"38815474",
   740 => x"81eb2e8c",
   741 => x"38805573",
   742 => x"752e0981",
   743 => x"0682f838",
   744 => x"80c5fb0b",
   745 => x"80f52d55",
   746 => x"748e3880",
   747 => x"c5fc0b80",
   748 => x"f52d5473",
   749 => x"822e8638",
   750 => x"80559a97",
   751 => x"0480c5fd",
   752 => x"0b80f52d",
   753 => x"7080cbf4",
   754 => x"0cff0580",
   755 => x"cbf80c80",
   756 => x"c5fe0b80",
   757 => x"f52d80c5",
   758 => x"ff0b80f5",
   759 => x"2d587605",
   760 => x"77828029",
   761 => x"057080cc",
   762 => x"840c80c6",
   763 => x"800b80f5",
   764 => x"2d7080cc",
   765 => x"980c80cb",
   766 => x"fc085957",
   767 => x"5876802e",
   768 => x"81b63888",
   769 => x"53be8c52",
   770 => x"80c6c251",
   771 => x"92ca2d80",
   772 => x"c2b80882",
   773 => x"823880cb",
   774 => x"f4087084",
   775 => x"2b80cc80",
   776 => x"0c7080cc",
   777 => x"940c80c6",
   778 => x"950b80f5",
   779 => x"2d80c694",
   780 => x"0b80f52d",
   781 => x"71828029",
   782 => x"0580c696",
   783 => x"0b80f52d",
   784 => x"70848080",
   785 => x"291280c6",
   786 => x"970b80f5",
   787 => x"2d708180",
   788 => x"0a291270",
   789 => x"80cc9c0c",
   790 => x"80cc9808",
   791 => x"712980cc",
   792 => x"84080570",
   793 => x"80cc880c",
   794 => x"80c69d0b",
   795 => x"80f52d80",
   796 => x"c69c0b80",
   797 => x"f52d7182",
   798 => x"80290580",
   799 => x"c69e0b80",
   800 => x"f52d7084",
   801 => x"80802912",
   802 => x"80c69f0b",
   803 => x"80f52d70",
   804 => x"982b81f0",
   805 => x"0a067205",
   806 => x"7080cc8c",
   807 => x"0cfe117e",
   808 => x"29770580",
   809 => x"cc900c52",
   810 => x"59524354",
   811 => x"5e515259",
   812 => x"525d5759",
   813 => x"579a9004",
   814 => x"80c6820b",
   815 => x"80f52d80",
   816 => x"c6810b80",
   817 => x"f52d7182",
   818 => x"80290570",
   819 => x"80cc800c",
   820 => x"70a02983",
   821 => x"ff057089",
   822 => x"2a7080cc",
   823 => x"940c80c6",
   824 => x"870b80f5",
   825 => x"2d80c686",
   826 => x"0b80f52d",
   827 => x"71828029",
   828 => x"057080cc",
   829 => x"9c0c7b71",
   830 => x"291e7080",
   831 => x"cc900c7d",
   832 => x"80cc8c0c",
   833 => x"730580cc",
   834 => x"880c555e",
   835 => x"51515555",
   836 => x"80519389",
   837 => x"2d815574",
   838 => x"80c2b80c",
   839 => x"02a8050d",
   840 => x"0402ec05",
   841 => x"0d767087",
   842 => x"2c7180ff",
   843 => x"06555654",
   844 => x"80cbfc08",
   845 => x"8a387388",
   846 => x"2c7481ff",
   847 => x"06545580",
   848 => x"c5f05280",
   849 => x"cc840815",
   850 => x"51a8812d",
   851 => x"80c2b808",
   852 => x"5480c2b8",
   853 => x"08802eb8",
   854 => x"3880cbfc",
   855 => x"08802e9a",
   856 => x"38728429",
   857 => x"80c5f005",
   858 => x"70085253",
   859 => x"a9a42d80",
   860 => x"c2b808f0",
   861 => x"0a06539b",
   862 => x"8e047210",
   863 => x"80c5f005",
   864 => x"7080e02d",
   865 => x"5253a9d5",
   866 => x"2d80c2b8",
   867 => x"08537254",
   868 => x"7380c2b8",
   869 => x"0c029405",
   870 => x"0d0402e0",
   871 => x"050d7970",
   872 => x"842c80cc",
   873 => x"a4080571",
   874 => x"8f065255",
   875 => x"53728a38",
   876 => x"80c5f052",
   877 => x"7351a881",
   878 => x"2d72a029",
   879 => x"80c5f005",
   880 => x"54807480",
   881 => x"f52d5653",
   882 => x"74732e83",
   883 => x"38815374",
   884 => x"81e52e81",
   885 => x"f4388170",
   886 => x"74065458",
   887 => x"72802e81",
   888 => x"e8388b14",
   889 => x"80f52d70",
   890 => x"832a7906",
   891 => x"5856769b",
   892 => x"3880c1e8",
   893 => x"08537289",
   894 => x"387280c9",
   895 => x"f00b81b7",
   896 => x"2d7680c1",
   897 => x"e80c7353",
   898 => x"9dcb0475",
   899 => x"8f2e0981",
   900 => x"0681b638",
   901 => x"749f068d",
   902 => x"2980c9e3",
   903 => x"11515381",
   904 => x"1480f52d",
   905 => x"73708105",
   906 => x"5581b72d",
   907 => x"831480f5",
   908 => x"2d737081",
   909 => x"055581b7",
   910 => x"2d851480",
   911 => x"f52d7370",
   912 => x"81055581",
   913 => x"b72d8714",
   914 => x"80f52d73",
   915 => x"70810555",
   916 => x"81b72d89",
   917 => x"1480f52d",
   918 => x"73708105",
   919 => x"5581b72d",
   920 => x"8e1480f5",
   921 => x"2d737081",
   922 => x"055581b7",
   923 => x"2d901480",
   924 => x"f52d7370",
   925 => x"81055581",
   926 => x"b72d9214",
   927 => x"80f52d73",
   928 => x"70810555",
   929 => x"81b72d94",
   930 => x"1480f52d",
   931 => x"73708105",
   932 => x"5581b72d",
   933 => x"961480f5",
   934 => x"2d737081",
   935 => x"055581b7",
   936 => x"2d981480",
   937 => x"f52d7370",
   938 => x"81055581",
   939 => x"b72d9c14",
   940 => x"80f52d73",
   941 => x"70810555",
   942 => x"81b72d9e",
   943 => x"1480f52d",
   944 => x"7381b72d",
   945 => x"7780c1e8",
   946 => x"0c805372",
   947 => x"80c2b80c",
   948 => x"02a0050d",
   949 => x"0402cc05",
   950 => x"0d7e605e",
   951 => x"5a800b80",
   952 => x"cca00880",
   953 => x"cca40859",
   954 => x"5c568058",
   955 => x"80cc8008",
   956 => x"782e81b8",
   957 => x"38778f06",
   958 => x"a0175754",
   959 => x"73913880",
   960 => x"c5f05276",
   961 => x"51811757",
   962 => x"a8812d80",
   963 => x"c5f05680",
   964 => x"7680f52d",
   965 => x"56547474",
   966 => x"2e833881",
   967 => x"547481e5",
   968 => x"2e80fd38",
   969 => x"81707506",
   970 => x"555c7380",
   971 => x"2e80f138",
   972 => x"8b1680f5",
   973 => x"2d980659",
   974 => x"7880e538",
   975 => x"8b537c52",
   976 => x"755192ca",
   977 => x"2d80c2b8",
   978 => x"0880d538",
   979 => x"9c160851",
   980 => x"a9a42d80",
   981 => x"c2b80884",
   982 => x"1b0c9a16",
   983 => x"80e02d51",
   984 => x"a9d52d80",
   985 => x"c2b80880",
   986 => x"c2b80888",
   987 => x"1c0c80c2",
   988 => x"b8085555",
   989 => x"80cbfc08",
   990 => x"802e9938",
   991 => x"941680e0",
   992 => x"2d51a9d5",
   993 => x"2d80c2b8",
   994 => x"08902b83",
   995 => x"fff00a06",
   996 => x"70165154",
   997 => x"73881b0c",
   998 => x"787a0c7b",
   999 => x"549fe804",
  1000 => x"81185880",
  1001 => x"cc800878",
  1002 => x"26feca38",
  1003 => x"80cbfc08",
  1004 => x"802eb338",
  1005 => x"7a519aa1",
  1006 => x"2d80c2b8",
  1007 => x"0880c2b8",
  1008 => x"0880ffff",
  1009 => x"fff80655",
  1010 => x"5b7380ff",
  1011 => x"fffff82e",
  1012 => x"953880c2",
  1013 => x"b808fe05",
  1014 => x"80cbf408",
  1015 => x"2980cc88",
  1016 => x"0805579d",
  1017 => x"ea048054",
  1018 => x"7380c2b8",
  1019 => x"0c02b405",
  1020 => x"0d0402f4",
  1021 => x"050d7470",
  1022 => x"08810571",
  1023 => x"0c700880",
  1024 => x"cbf80806",
  1025 => x"5353718f",
  1026 => x"38881308",
  1027 => x"519aa12d",
  1028 => x"80c2b808",
  1029 => x"88140c81",
  1030 => x"0b80c2b8",
  1031 => x"0c028c05",
  1032 => x"0d0402f0",
  1033 => x"050d7588",
  1034 => x"1108fe05",
  1035 => x"80cbf408",
  1036 => x"2980cc88",
  1037 => x"08117208",
  1038 => x"80cbf808",
  1039 => x"06057955",
  1040 => x"535454a8",
  1041 => x"812d0290",
  1042 => x"050d0402",
  1043 => x"f0050d75",
  1044 => x"881108fe",
  1045 => x"0580cbf4",
  1046 => x"082980cc",
  1047 => x"88081172",
  1048 => x"0880cbf8",
  1049 => x"08060579",
  1050 => x"55535454",
  1051 => x"a6bf2d02",
  1052 => x"90050d04",
  1053 => x"02f4050d",
  1054 => x"d45281ff",
  1055 => x"720c7108",
  1056 => x"5381ff72",
  1057 => x"0c72882b",
  1058 => x"83fe8006",
  1059 => x"72087081",
  1060 => x"ff065152",
  1061 => x"5381ff72",
  1062 => x"0c727107",
  1063 => x"882b7208",
  1064 => x"7081ff06",
  1065 => x"51525381",
  1066 => x"ff720c72",
  1067 => x"7107882b",
  1068 => x"72087081",
  1069 => x"ff067207",
  1070 => x"80c2b80c",
  1071 => x"5253028c",
  1072 => x"050d0402",
  1073 => x"f4050d74",
  1074 => x"767181ff",
  1075 => x"06d40c53",
  1076 => x"5380ccac",
  1077 => x"08853871",
  1078 => x"892b5271",
  1079 => x"982ad40c",
  1080 => x"71902a70",
  1081 => x"81ff06d4",
  1082 => x"0c517188",
  1083 => x"2a7081ff",
  1084 => x"06d40c51",
  1085 => x"7181ff06",
  1086 => x"d40c7290",
  1087 => x"2a7081ff",
  1088 => x"06d40c51",
  1089 => x"d4087081",
  1090 => x"ff065151",
  1091 => x"82b8bf52",
  1092 => x"7081ff2e",
  1093 => x"09810694",
  1094 => x"3881ff0b",
  1095 => x"d40cd408",
  1096 => x"7081ff06",
  1097 => x"ff145451",
  1098 => x"5171e538",
  1099 => x"7080c2b8",
  1100 => x"0c028c05",
  1101 => x"0d0402fc",
  1102 => x"050d81c7",
  1103 => x"5181ff0b",
  1104 => x"d40cff11",
  1105 => x"51708025",
  1106 => x"f4380284",
  1107 => x"050d0402",
  1108 => x"f0050da2",
  1109 => x"b62d8fcf",
  1110 => x"53805287",
  1111 => x"fc80f751",
  1112 => x"a1c32d80",
  1113 => x"c2b80854",
  1114 => x"80c2b808",
  1115 => x"812e0981",
  1116 => x"06a43881",
  1117 => x"ff0bd40c",
  1118 => x"820a5284",
  1119 => x"9c80e951",
  1120 => x"a1c32d80",
  1121 => x"c2b8088b",
  1122 => x"3881ff0b",
  1123 => x"d40c7353",
  1124 => x"a39d04a2",
  1125 => x"b62dff13",
  1126 => x"5372ffbd",
  1127 => x"387280c2",
  1128 => x"b80c0290",
  1129 => x"050d0402",
  1130 => x"f4050d81",
  1131 => x"ff0bd40c",
  1132 => x"93538052",
  1133 => x"87fc80c1",
  1134 => x"51a1c32d",
  1135 => x"80c2b808",
  1136 => x"8b3881ff",
  1137 => x"0bd40c81",
  1138 => x"53a3d504",
  1139 => x"a2b62dff",
  1140 => x"135372de",
  1141 => x"387280c2",
  1142 => x"b80c028c",
  1143 => x"050d0402",
  1144 => x"f0050da2",
  1145 => x"b62d83aa",
  1146 => x"52849c80",
  1147 => x"c851a1c3",
  1148 => x"2d80c2b8",
  1149 => x"08812e09",
  1150 => x"81069338",
  1151 => x"a0f42d80",
  1152 => x"c2b80883",
  1153 => x"ffff0653",
  1154 => x"7283aa2e",
  1155 => x"9738a3a7",
  1156 => x"2da49f04",
  1157 => x"8154a587",
  1158 => x"04beb851",
  1159 => x"86922d80",
  1160 => x"54a58704",
  1161 => x"81ff0bd4",
  1162 => x"0cb153a2",
  1163 => x"cf2d80c2",
  1164 => x"b808802e",
  1165 => x"80c23880",
  1166 => x"5287fc80",
  1167 => x"fa51a1c3",
  1168 => x"2d80c2b8",
  1169 => x"08b23881",
  1170 => x"ff0bd40c",
  1171 => x"d4085381",
  1172 => x"ff0bd40c",
  1173 => x"81ff0bd4",
  1174 => x"0c81ff0b",
  1175 => x"d40c81ff",
  1176 => x"0bd40c72",
  1177 => x"862a7081",
  1178 => x"0680c2b8",
  1179 => x"08565153",
  1180 => x"72802e93",
  1181 => x"38a49404",
  1182 => x"72822eff",
  1183 => x"9c38ff13",
  1184 => x"5372ffa7",
  1185 => x"38725473",
  1186 => x"80c2b80c",
  1187 => x"0290050d",
  1188 => x"0402f005",
  1189 => x"0d810b80",
  1190 => x"ccac0c84",
  1191 => x"54d00870",
  1192 => x"8f2a7081",
  1193 => x"06515153",
  1194 => x"72f33872",
  1195 => x"d00ca2b6",
  1196 => x"2dbec851",
  1197 => x"86922dd0",
  1198 => x"08708f2a",
  1199 => x"70810651",
  1200 => x"515372f3",
  1201 => x"38810bd0",
  1202 => x"0cb15380",
  1203 => x"5284d480",
  1204 => x"c051a1c3",
  1205 => x"2d80c2b8",
  1206 => x"08812ea1",
  1207 => x"3872822e",
  1208 => x"0981068c",
  1209 => x"38bed451",
  1210 => x"86922d80",
  1211 => x"53a6b504",
  1212 => x"ff135372",
  1213 => x"d638ff14",
  1214 => x"5473ffa1",
  1215 => x"38a3df2d",
  1216 => x"80c2b808",
  1217 => x"80ccac0c",
  1218 => x"80c2b808",
  1219 => x"8b388152",
  1220 => x"87fc80d0",
  1221 => x"51a1c32d",
  1222 => x"81ff0bd4",
  1223 => x"0cd00870",
  1224 => x"8f2a7081",
  1225 => x"06515153",
  1226 => x"72f33872",
  1227 => x"d00c81ff",
  1228 => x"0bd40c81",
  1229 => x"537280c2",
  1230 => x"b80c0290",
  1231 => x"050d0402",
  1232 => x"e8050d78",
  1233 => x"5681ff0b",
  1234 => x"d40cd008",
  1235 => x"708f2a70",
  1236 => x"81065151",
  1237 => x"5372f338",
  1238 => x"82810bd0",
  1239 => x"0c81ff0b",
  1240 => x"d40c7752",
  1241 => x"87fc80d8",
  1242 => x"51a1c32d",
  1243 => x"80c2b808",
  1244 => x"802e8c38",
  1245 => x"beec5186",
  1246 => x"922d8153",
  1247 => x"a7f70481",
  1248 => x"ff0bd40c",
  1249 => x"81fe0bd4",
  1250 => x"0c80ff55",
  1251 => x"75708405",
  1252 => x"57087098",
  1253 => x"2ad40c70",
  1254 => x"902c7081",
  1255 => x"ff06d40c",
  1256 => x"5470882c",
  1257 => x"7081ff06",
  1258 => x"d40c5470",
  1259 => x"81ff06d4",
  1260 => x"0c54ff15",
  1261 => x"55748025",
  1262 => x"d33881ff",
  1263 => x"0bd40c81",
  1264 => x"ff0bd40c",
  1265 => x"81ff0bd4",
  1266 => x"0c868da0",
  1267 => x"5481ff0b",
  1268 => x"d40cd408",
  1269 => x"81ff0655",
  1270 => x"748738ff",
  1271 => x"145473ed",
  1272 => x"3881ff0b",
  1273 => x"d40cd008",
  1274 => x"708f2a70",
  1275 => x"81065151",
  1276 => x"5372f338",
  1277 => x"72d00c72",
  1278 => x"80c2b80c",
  1279 => x"0298050d",
  1280 => x"0402e805",
  1281 => x"0d785580",
  1282 => x"5681ff0b",
  1283 => x"d40cd008",
  1284 => x"708f2a70",
  1285 => x"81065151",
  1286 => x"5372f338",
  1287 => x"82810bd0",
  1288 => x"0c81ff0b",
  1289 => x"d40c7752",
  1290 => x"87fc80d1",
  1291 => x"51a1c32d",
  1292 => x"80dbc6df",
  1293 => x"5480c2b8",
  1294 => x"08802e8a",
  1295 => x"38befc51",
  1296 => x"86922da9",
  1297 => x"9a0481ff",
  1298 => x"0bd40cd4",
  1299 => x"087081ff",
  1300 => x"06515372",
  1301 => x"81fe2e09",
  1302 => x"81069e38",
  1303 => x"80ff53a0",
  1304 => x"f42d80c2",
  1305 => x"b8087570",
  1306 => x"8405570c",
  1307 => x"ff135372",
  1308 => x"8025ec38",
  1309 => x"8156a8ff",
  1310 => x"04ff1454",
  1311 => x"73c83881",
  1312 => x"ff0bd40c",
  1313 => x"81ff0bd4",
  1314 => x"0cd00870",
  1315 => x"8f2a7081",
  1316 => x"06515153",
  1317 => x"72f33872",
  1318 => x"d00c7580",
  1319 => x"c2b80c02",
  1320 => x"98050d04",
  1321 => x"02f4050d",
  1322 => x"7470882a",
  1323 => x"83fe8006",
  1324 => x"7072982a",
  1325 => x"0772882b",
  1326 => x"87fc8080",
  1327 => x"0673982b",
  1328 => x"81f00a06",
  1329 => x"71730707",
  1330 => x"80c2b80c",
  1331 => x"56515351",
  1332 => x"028c050d",
  1333 => x"0402f805",
  1334 => x"0d028e05",
  1335 => x"80f52d74",
  1336 => x"882b0770",
  1337 => x"83ffff06",
  1338 => x"80c2b80c",
  1339 => x"51028805",
  1340 => x"0d0402fc",
  1341 => x"050d7251",
  1342 => x"80710c80",
  1343 => x"0b84120c",
  1344 => x"0284050d",
  1345 => x"0402f005",
  1346 => x"0d757008",
  1347 => x"84120853",
  1348 => x"5353ff54",
  1349 => x"71712ea8",
  1350 => x"38addc2d",
  1351 => x"84130870",
  1352 => x"84291488",
  1353 => x"11700870",
  1354 => x"81ff0684",
  1355 => x"18088111",
  1356 => x"8706841a",
  1357 => x"0c535155",
  1358 => x"515151ad",
  1359 => x"d62d7154",
  1360 => x"7380c2b8",
  1361 => x"0c029005",
  1362 => x"0d0402f8",
  1363 => x"050daddc",
  1364 => x"2de00870",
  1365 => x"8b2a7081",
  1366 => x"06515252",
  1367 => x"70802ea1",
  1368 => x"3880ccb0",
  1369 => x"08708429",
  1370 => x"80ccb805",
  1371 => x"7381ff06",
  1372 => x"710c5151",
  1373 => x"80ccb008",
  1374 => x"81118706",
  1375 => x"80ccb00c",
  1376 => x"51800b80",
  1377 => x"ccd80cad",
  1378 => x"ce2dadd6",
  1379 => x"2d028805",
  1380 => x"0d0402fc",
  1381 => x"050daddc",
  1382 => x"2d810b80",
  1383 => x"ccd80cad",
  1384 => x"d62d80cc",
  1385 => x"d8085170",
  1386 => x"f9380284",
  1387 => x"050d0402",
  1388 => x"fc050d80",
  1389 => x"ccb051a9",
  1390 => x"f22daaca",
  1391 => x"51adca2d",
  1392 => x"acf12d02",
  1393 => x"84050d04",
  1394 => x"02f4050d",
  1395 => x"acd60480",
  1396 => x"c2b80881",
  1397 => x"f02e0981",
  1398 => x"068a3881",
  1399 => x"0b80c2ac",
  1400 => x"0cacd604",
  1401 => x"80c2b808",
  1402 => x"81e02e09",
  1403 => x"81068a38",
  1404 => x"810b80c2",
  1405 => x"b00cacd6",
  1406 => x"0480c2b8",
  1407 => x"085280c2",
  1408 => x"b008802e",
  1409 => x"893880c2",
  1410 => x"b8088180",
  1411 => x"05527184",
  1412 => x"2c728f06",
  1413 => x"535380c2",
  1414 => x"ac08802e",
  1415 => x"9a387284",
  1416 => x"2980c1ec",
  1417 => x"05721381",
  1418 => x"712b7009",
  1419 => x"73080673",
  1420 => x"0c515353",
  1421 => x"acca0472",
  1422 => x"842980c1",
  1423 => x"ec057213",
  1424 => x"83712b72",
  1425 => x"0807720c",
  1426 => x"5353800b",
  1427 => x"80c2b00c",
  1428 => x"800b80c2",
  1429 => x"ac0c80cc",
  1430 => x"b051aa85",
  1431 => x"2d80c2b8",
  1432 => x"08ff24fe",
  1433 => x"ea38800b",
  1434 => x"80c2b80c",
  1435 => x"028c050d",
  1436 => x"0402f805",
  1437 => x"0d80c1ec",
  1438 => x"528f5180",
  1439 => x"72708405",
  1440 => x"540cff11",
  1441 => x"51708025",
  1442 => x"f2380288",
  1443 => x"050d0402",
  1444 => x"f0050d75",
  1445 => x"51addc2d",
  1446 => x"70822cfc",
  1447 => x"0680c1ec",
  1448 => x"1172109e",
  1449 => x"06710870",
  1450 => x"722a7083",
  1451 => x"0682742b",
  1452 => x"70097406",
  1453 => x"760c5451",
  1454 => x"56575351",
  1455 => x"53add62d",
  1456 => x"7180c2b8",
  1457 => x"0c029005",
  1458 => x"0d047198",
  1459 => x"0c04ffb0",
  1460 => x"0880c2b8",
  1461 => x"0c04810b",
  1462 => x"ffb00c04",
  1463 => x"800bffb0",
  1464 => x"0c0402fc",
  1465 => x"050d810b",
  1466 => x"80c2b40c",
  1467 => x"81518581",
  1468 => x"2d028405",
  1469 => x"0d0402fc",
  1470 => x"050d800b",
  1471 => x"80c2b40c",
  1472 => x"80518581",
  1473 => x"2d028405",
  1474 => x"0d0402ec",
  1475 => x"050d7654",
  1476 => x"8052870b",
  1477 => x"881580f5",
  1478 => x"2d565374",
  1479 => x"72248338",
  1480 => x"a0537251",
  1481 => x"82f82d81",
  1482 => x"128b1580",
  1483 => x"f52d5452",
  1484 => x"727225de",
  1485 => x"38029405",
  1486 => x"0d0402f0",
  1487 => x"050d80cc",
  1488 => x"e8085481",
  1489 => x"f92d800b",
  1490 => x"80ccec0c",
  1491 => x"7308802e",
  1492 => x"81863882",
  1493 => x"0b80c2cc",
  1494 => x"0c80ccec",
  1495 => x"088f0680",
  1496 => x"c2c80c73",
  1497 => x"08527183",
  1498 => x"2e963871",
  1499 => x"83268938",
  1500 => x"71812eaf",
  1501 => x"38afc104",
  1502 => x"71852e9f",
  1503 => x"38afc104",
  1504 => x"881480f5",
  1505 => x"2d841508",
  1506 => x"bf8c5354",
  1507 => x"5286922d",
  1508 => x"71842913",
  1509 => x"70085252",
  1510 => x"afc50473",
  1511 => x"51ae8a2d",
  1512 => x"afc10480",
  1513 => x"ccdc0888",
  1514 => x"15082c70",
  1515 => x"81065152",
  1516 => x"71802e87",
  1517 => x"38bf9051",
  1518 => x"afbe04bf",
  1519 => x"94518692",
  1520 => x"2d841408",
  1521 => x"5186922d",
  1522 => x"80ccec08",
  1523 => x"810580cc",
  1524 => x"ec0c8c14",
  1525 => x"54aecc04",
  1526 => x"0290050d",
  1527 => x"047180cc",
  1528 => x"e80caeba",
  1529 => x"2d80ccec",
  1530 => x"08ff0580",
  1531 => x"ccf00c04",
  1532 => x"7180ccf4",
  1533 => x"0c0402e8",
  1534 => x"050d80cc",
  1535 => x"e80880cc",
  1536 => x"f4085755",
  1537 => x"80f851ad",
  1538 => x"8f2d80c2",
  1539 => x"b808812a",
  1540 => x"70810651",
  1541 => x"52719c38",
  1542 => x"8751ad8f",
  1543 => x"2d80c2b8",
  1544 => x"08812a70",
  1545 => x"81065152",
  1546 => x"71802eb5",
  1547 => x"38b0b304",
  1548 => x"abc82d87",
  1549 => x"51ad8f2d",
  1550 => x"80c2b808",
  1551 => x"f338b0c4",
  1552 => x"04abc82d",
  1553 => x"80f851ad",
  1554 => x"8f2d80c2",
  1555 => x"b808f238",
  1556 => x"80c2b408",
  1557 => x"81327080",
  1558 => x"c2b40c70",
  1559 => x"52528581",
  1560 => x"2d800b80",
  1561 => x"cce00c80",
  1562 => x"0b80cce4",
  1563 => x"0c80c2b4",
  1564 => x"08838d38",
  1565 => x"80da51ad",
  1566 => x"8f2d80c2",
  1567 => x"b808802e",
  1568 => x"8c3880cc",
  1569 => x"e0088180",
  1570 => x"0780cce0",
  1571 => x"0c80d951",
  1572 => x"ad8f2d80",
  1573 => x"c2b80880",
  1574 => x"2e8c3880",
  1575 => x"cce00880",
  1576 => x"c00780cc",
  1577 => x"e00c8194",
  1578 => x"51ad8f2d",
  1579 => x"80c2b808",
  1580 => x"802e8b38",
  1581 => x"80cce008",
  1582 => x"900780cc",
  1583 => x"e00c8191",
  1584 => x"51ad8f2d",
  1585 => x"80c2b808",
  1586 => x"802e8b38",
  1587 => x"80cce008",
  1588 => x"a00780cc",
  1589 => x"e00c81f5",
  1590 => x"51ad8f2d",
  1591 => x"80c2b808",
  1592 => x"802e8b38",
  1593 => x"80cce008",
  1594 => x"810780cc",
  1595 => x"e00c81f2",
  1596 => x"51ad8f2d",
  1597 => x"80c2b808",
  1598 => x"802e8b38",
  1599 => x"80cce008",
  1600 => x"820780cc",
  1601 => x"e00c81eb",
  1602 => x"51ad8f2d",
  1603 => x"80c2b808",
  1604 => x"802e8b38",
  1605 => x"80cce008",
  1606 => x"840780cc",
  1607 => x"e00c81f4",
  1608 => x"51ad8f2d",
  1609 => x"80c2b808",
  1610 => x"802e8b38",
  1611 => x"80cce008",
  1612 => x"880780cc",
  1613 => x"e00c80d8",
  1614 => x"51ad8f2d",
  1615 => x"80c2b808",
  1616 => x"802e8c38",
  1617 => x"80cce408",
  1618 => x"81800780",
  1619 => x"cce40c92",
  1620 => x"51ad8f2d",
  1621 => x"80c2b808",
  1622 => x"802e8c38",
  1623 => x"80cce408",
  1624 => x"80c00780",
  1625 => x"cce40c94",
  1626 => x"51ad8f2d",
  1627 => x"80c2b808",
  1628 => x"802e8b38",
  1629 => x"80cce408",
  1630 => x"900780cc",
  1631 => x"e40c9151",
  1632 => x"ad8f2d80",
  1633 => x"c2b80880",
  1634 => x"2e8b3880",
  1635 => x"cce408a0",
  1636 => x"0780cce4",
  1637 => x"0c9d51ad",
  1638 => x"8f2d80c2",
  1639 => x"b808802e",
  1640 => x"8b3880cc",
  1641 => x"e4088107",
  1642 => x"80cce40c",
  1643 => x"9b51ad8f",
  1644 => x"2d80c2b8",
  1645 => x"08802e8b",
  1646 => x"3880cce4",
  1647 => x"08820780",
  1648 => x"cce40c9c",
  1649 => x"51ad8f2d",
  1650 => x"80c2b808",
  1651 => x"802e8b38",
  1652 => x"80cce408",
  1653 => x"840780cc",
  1654 => x"e40ca351",
  1655 => x"ad8f2d80",
  1656 => x"c2b80880",
  1657 => x"2e8b3880",
  1658 => x"cce40888",
  1659 => x"0780cce4",
  1660 => x"0c81fd51",
  1661 => x"ad8f2d81",
  1662 => x"fa51ad8f",
  1663 => x"2db9d504",
  1664 => x"81f551ad",
  1665 => x"8f2d80c2",
  1666 => x"b808812a",
  1667 => x"70810651",
  1668 => x"5271802e",
  1669 => x"b33880cc",
  1670 => x"f0085271",
  1671 => x"802e8a38",
  1672 => x"ff1280cc",
  1673 => x"f00cb4c8",
  1674 => x"0480ccec",
  1675 => x"081080cc",
  1676 => x"ec080570",
  1677 => x"84291651",
  1678 => x"52881208",
  1679 => x"802e8938",
  1680 => x"ff518812",
  1681 => x"0852712d",
  1682 => x"81f251ad",
  1683 => x"8f2d80c2",
  1684 => x"b808812a",
  1685 => x"70810651",
  1686 => x"5271802e",
  1687 => x"b43880cc",
  1688 => x"ec08ff11",
  1689 => x"80ccf008",
  1690 => x"56535373",
  1691 => x"72258a38",
  1692 => x"811480cc",
  1693 => x"f00cb591",
  1694 => x"04721013",
  1695 => x"70842916",
  1696 => x"51528812",
  1697 => x"08802e89",
  1698 => x"38fe5188",
  1699 => x"12085271",
  1700 => x"2d81fd51",
  1701 => x"ad8f2d80",
  1702 => x"c2b80881",
  1703 => x"2a708106",
  1704 => x"51527180",
  1705 => x"2eb13880",
  1706 => x"ccf00880",
  1707 => x"2e8a3880",
  1708 => x"0b80ccf0",
  1709 => x"0cb5d704",
  1710 => x"80ccec08",
  1711 => x"1080ccec",
  1712 => x"08057084",
  1713 => x"29165152",
  1714 => x"88120880",
  1715 => x"2e8938fd",
  1716 => x"51881208",
  1717 => x"52712d81",
  1718 => x"fa51ad8f",
  1719 => x"2d80c2b8",
  1720 => x"08812a70",
  1721 => x"81065152",
  1722 => x"71802eb1",
  1723 => x"3880ccec",
  1724 => x"08ff1154",
  1725 => x"5280ccf0",
  1726 => x"08732589",
  1727 => x"387280cc",
  1728 => x"f00cb69d",
  1729 => x"04711012",
  1730 => x"70842916",
  1731 => x"51528812",
  1732 => x"08802e89",
  1733 => x"38fc5188",
  1734 => x"12085271",
  1735 => x"2d80ccf0",
  1736 => x"08705354",
  1737 => x"73802e8a",
  1738 => x"388c15ff",
  1739 => x"155555b6",
  1740 => x"a404820b",
  1741 => x"80c2cc0c",
  1742 => x"718f0680",
  1743 => x"c2c80c81",
  1744 => x"eb51ad8f",
  1745 => x"2d80c2b8",
  1746 => x"08812a70",
  1747 => x"81065152",
  1748 => x"71802ead",
  1749 => x"38740885",
  1750 => x"2e098106",
  1751 => x"a4388815",
  1752 => x"80f52dff",
  1753 => x"05527188",
  1754 => x"1681b72d",
  1755 => x"71982b52",
  1756 => x"71802588",
  1757 => x"38800b88",
  1758 => x"1681b72d",
  1759 => x"7451ae8a",
  1760 => x"2d81f451",
  1761 => x"ad8f2d80",
  1762 => x"c2b80881",
  1763 => x"2a708106",
  1764 => x"51527180",
  1765 => x"2eb33874",
  1766 => x"08852e09",
  1767 => x"8106aa38",
  1768 => x"881580f5",
  1769 => x"2d810552",
  1770 => x"71881681",
  1771 => x"b72d7181",
  1772 => x"ff068b16",
  1773 => x"80f52d54",
  1774 => x"52727227",
  1775 => x"87387288",
  1776 => x"1681b72d",
  1777 => x"7451ae8a",
  1778 => x"2d80da51",
  1779 => x"ad8f2d80",
  1780 => x"c2b80881",
  1781 => x"2a708106",
  1782 => x"51527180",
  1783 => x"2e81ad38",
  1784 => x"80cce808",
  1785 => x"80ccf008",
  1786 => x"55537380",
  1787 => x"2e8a388c",
  1788 => x"13ff1555",
  1789 => x"53b7ea04",
  1790 => x"72085271",
  1791 => x"822ea638",
  1792 => x"71822689",
  1793 => x"3871812e",
  1794 => x"aa38b98c",
  1795 => x"0471832e",
  1796 => x"b4387184",
  1797 => x"2e098106",
  1798 => x"80f23888",
  1799 => x"130851af",
  1800 => x"dd2db98c",
  1801 => x"0480ccf0",
  1802 => x"08518813",
  1803 => x"0852712d",
  1804 => x"b98c0481",
  1805 => x"0b881408",
  1806 => x"2b80ccdc",
  1807 => x"083280cc",
  1808 => x"dc0cb8e0",
  1809 => x"04881380",
  1810 => x"f52d8105",
  1811 => x"8b1480f5",
  1812 => x"2d535471",
  1813 => x"74248338",
  1814 => x"80547388",
  1815 => x"1481b72d",
  1816 => x"aeba2db9",
  1817 => x"8c047508",
  1818 => x"802ea438",
  1819 => x"750851ad",
  1820 => x"8f2d80c2",
  1821 => x"b8088106",
  1822 => x"5271802e",
  1823 => x"8c3880cc",
  1824 => x"f0085184",
  1825 => x"16085271",
  1826 => x"2d881656",
  1827 => x"75d83880",
  1828 => x"54800b80",
  1829 => x"c2cc0c73",
  1830 => x"8f0680c2",
  1831 => x"c80ca052",
  1832 => x"7380ccf0",
  1833 => x"082e0981",
  1834 => x"06993880",
  1835 => x"ccec08ff",
  1836 => x"05743270",
  1837 => x"09810570",
  1838 => x"72079f2a",
  1839 => x"91713151",
  1840 => x"51535371",
  1841 => x"5182f82d",
  1842 => x"8114548e",
  1843 => x"7425c238",
  1844 => x"80c2b408",
  1845 => x"527180c2",
  1846 => x"b80c0298",
  1847 => x"050d0402",
  1848 => x"f0050d75",
  1849 => x"53875472",
  1850 => x"9c2ab005",
  1851 => x"52b97227",
  1852 => x"84388712",
  1853 => x"52715182",
  1854 => x"f82d7284",
  1855 => x"2bff1555",
  1856 => x"53738025",
  1857 => x"e2380290",
  1858 => x"050d0402",
  1859 => x"d4050d81",
  1860 => x"5481f92d",
  1861 => x"bbf104ff",
  1862 => x"145473a0",
  1863 => x"3887e854",
  1864 => x"ff707172",
  1865 => x"80c2b808",
  1866 => x"80c2b808",
  1867 => x"80c2b808",
  1868 => x"80c2b808",
  1869 => x"5c5c5c5c",
  1870 => x"5c5c5c53",
  1871 => x"80c2b808",
  1872 => x"80c2cc0c",
  1873 => x"80c2b808",
  1874 => x"80c2c80c",
  1875 => x"f4800870",
  1876 => x"7c067872",
  1877 => x"07595c51",
  1878 => x"b9df2da0",
  1879 => x"5182f82d",
  1880 => x"7a51b9df",
  1881 => x"2da05182",
  1882 => x"f82d7651",
  1883 => x"b9df2d8a",
  1884 => x"5182f82d",
  1885 => x"f4840870",
  1886 => x"74067972",
  1887 => x"075a5451",
  1888 => x"b9df2da0",
  1889 => x"5182f82d",
  1890 => x"7251b9df",
  1891 => x"2da05182",
  1892 => x"f82d7751",
  1893 => x"b9df2d8a",
  1894 => x"5182f82d",
  1895 => x"f4880870",
  1896 => x"7a067672",
  1897 => x"07575a51",
  1898 => x"b9df2da0",
  1899 => x"5182f82d",
  1900 => x"7851b9df",
  1901 => x"2da05182",
  1902 => x"f82d7451",
  1903 => x"b9df2d8a",
  1904 => x"5182f82d",
  1905 => x"f48c0870",
  1906 => x"7b067772",
  1907 => x"07725458",
  1908 => x"5b52b9df",
  1909 => x"2da05182",
  1910 => x"f82d7951",
  1911 => x"b9df2da0",
  1912 => x"5182f82d",
  1913 => x"7551b9df",
  1914 => x"2d8a5182",
  1915 => x"f82dabc8",
  1916 => x"2d80f651",
  1917 => x"ad8f2d80",
  1918 => x"c2b80880",
  1919 => x"2efe9838",
  1920 => x"aeba2d71",
  1921 => x"80c2b80c",
  1922 => x"02ac050d",
  1923 => x"04000000",
  1924 => x"00ffffff",
  1925 => x"ff00ffff",
  1926 => x"ffff00ff",
  1927 => x"ffffff00",
  1928 => x"52657365",
  1929 => x"74000000",
  1930 => x"53617665",
  1931 => x"20736574",
  1932 => x"74696e67",
  1933 => x"73000000",
  1934 => x"5363616e",
  1935 => x"6c696e65",
  1936 => x"73000000",
  1937 => x"4c6f6164",
  1938 => x"20524f4d",
  1939 => x"20100000",
  1940 => x"44656275",
  1941 => x"67201000",
  1942 => x"45786974",
  1943 => x"00000000",
  1944 => x"50432045",
  1945 => x"6e67696e",
  1946 => x"65206d6f",
  1947 => x"64650000",
  1948 => x"54757262",
  1949 => x"6f677261",
  1950 => x"66782031",
  1951 => x"36206d6f",
  1952 => x"64650000",
  1953 => x"56474120",
  1954 => x"2d203331",
  1955 => x"4b487a2c",
  1956 => x"20363048",
  1957 => x"7a000000",
  1958 => x"5456202d",
  1959 => x"20343830",
  1960 => x"692c2036",
  1961 => x"30487a00",
  1962 => x"4261636b",
  1963 => x"00000000",
  1964 => x"46504741",
  1965 => x"50434520",
  1966 => x"43464700",
  1967 => x"496e6974",
  1968 => x"69616c69",
  1969 => x"7a696e67",
  1970 => x"20534420",
  1971 => x"63617264",
  1972 => x"0a000000",
  1973 => x"424f4f54",
  1974 => x"20202020",
  1975 => x"50434500",
  1976 => x"43617264",
  1977 => x"20696e69",
  1978 => x"74206661",
  1979 => x"696c6564",
  1980 => x"0a000000",
  1981 => x"4d425220",
  1982 => x"6661696c",
  1983 => x"0a000000",
  1984 => x"46415431",
  1985 => x"36202020",
  1986 => x"00000000",
  1987 => x"46415433",
  1988 => x"32202020",
  1989 => x"00000000",
  1990 => x"4e6f2070",
  1991 => x"61727469",
  1992 => x"74696f6e",
  1993 => x"20736967",
  1994 => x"0a000000",
  1995 => x"42616420",
  1996 => x"70617274",
  1997 => x"0a000000",
  1998 => x"53444843",
  1999 => x"20657272",
  2000 => x"6f72210a",
  2001 => x"00000000",
  2002 => x"53442069",
  2003 => x"6e69742e",
  2004 => x"2e2e0a00",
  2005 => x"53442063",
  2006 => x"61726420",
  2007 => x"72657365",
  2008 => x"74206661",
  2009 => x"696c6564",
  2010 => x"210a0000",
  2011 => x"57726974",
  2012 => x"65206661",
  2013 => x"696c6564",
  2014 => x"0a000000",
  2015 => x"52656164",
  2016 => x"20666169",
  2017 => x"6c65640a",
  2018 => x"00000000",
  2019 => x"16200000",
  2020 => x"14200000",
  2021 => x"15200000",
  2022 => x"00000002",
  2023 => x"00000002",
  2024 => x"00001e20",
  2025 => x"000004f4",
  2026 => x"00000002",
  2027 => x"00001e28",
  2028 => x"000003a2",
  2029 => x"00000003",
  2030 => x"00002010",
  2031 => x"00000002",
  2032 => x"00000001",
  2033 => x"00001e38",
  2034 => x"00000001",
  2035 => x"00000003",
  2036 => x"00002008",
  2037 => x"00000002",
  2038 => x"00000002",
  2039 => x"00001e44",
  2040 => x"000007e3",
  2041 => x"00000002",
  2042 => x"00001e50",
  2043 => x"00001d0b",
  2044 => x"00000002",
  2045 => x"00001e58",
  2046 => x"000016f6",
  2047 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

