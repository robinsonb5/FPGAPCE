-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb2",
     9 => x"fc080b0b",
    10 => x"0bb38008",
    11 => x"0b0b0bb3",
    12 => x"84080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b3840c0b",
    16 => x"0b0bb380",
    17 => x"0c0b0b0b",
    18 => x"b2fc0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bace8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b2fc70b9",
    57 => x"e8278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8ccf0402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b38c0c9f",
    65 => x"0bb3900c",
    66 => x"a0717081",
    67 => x"055334b3",
    68 => x"9008ff05",
    69 => x"b3900cb3",
    70 => x"90088025",
    71 => x"eb38b38c",
    72 => x"08ff05b3",
    73 => x"8c0cb38c",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb38c",
    94 => x"08258f38",
    95 => x"82b22db3",
    96 => x"8c08ff05",
    97 => x"b38c0c82",
    98 => x"f404b38c",
    99 => x"08b39008",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b38c08",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b3",
   108 => x"90088105",
   109 => x"b3900cb3",
   110 => x"9008519f",
   111 => x"7125e238",
   112 => x"800bb390",
   113 => x"0cb38c08",
   114 => x"8105b38c",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b3900881",
   120 => x"05b3900c",
   121 => x"b39008a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b3900cb3",
   125 => x"8c088105",
   126 => x"b38c0c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb3",
   155 => x"940cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb394",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b3940884",
   167 => x"07b3940c",
   168 => x"5573842b",
   169 => x"87e87125",
   170 => x"83713170",
   171 => x"0b0b0bb0",
   172 => x"840c8171",
   173 => x"2bf6880c",
   174 => x"fea413ff",
   175 => x"122c7888",
   176 => x"29ff9405",
   177 => x"70812cb3",
   178 => x"94085258",
   179 => x"52555152",
   180 => x"5476802e",
   181 => x"85387081",
   182 => x"075170f6",
   183 => x"940c7109",
   184 => x"8105f680",
   185 => x"0c720981",
   186 => x"05f6840c",
   187 => x"0294050d",
   188 => x"0402f405",
   189 => x"0d745372",
   190 => x"70810554",
   191 => x"80f52d52",
   192 => x"71802e89",
   193 => x"38715182",
   194 => x"ee2d85f7",
   195 => x"04028c05",
   196 => x"0d0402f4",
   197 => x"050d7470",
   198 => x"8206b9d8",
   199 => x"0cb0a071",
   200 => x"81065454",
   201 => x"51718814",
   202 => x"81b72d70",
   203 => x"822a7081",
   204 => x"06515170",
   205 => x"941481b7",
   206 => x"2d70b2fc",
   207 => x"0c028c05",
   208 => x"0d0402f4",
   209 => x"050dae80",
   210 => x"52b39c51",
   211 => x"95df2db2",
   212 => x"fc08802e",
   213 => x"9538b4f8",
   214 => x"52b39c51",
   215 => x"98952db4",
   216 => x"f80870fe",
   217 => x"c00c5186",
   218 => x"922d028c",
   219 => x"050d0402",
   220 => x"f8050db9",
   221 => x"d8088206",
   222 => x"b0a80b80",
   223 => x"f52d5252",
   224 => x"70802e85",
   225 => x"38718107",
   226 => x"52b0b40b",
   227 => x"80f52d51",
   228 => x"70802e85",
   229 => x"38718407",
   230 => x"5271b2fc",
   231 => x"0c028805",
   232 => x"0d0402f0",
   233 => x"050d86ef",
   234 => x"2db2fc08",
   235 => x"ae8053b3",
   236 => x"9c525395",
   237 => x"df2db2fc",
   238 => x"08802ea3",
   239 => x"3872b4f8",
   240 => x"0cb4fc54",
   241 => x"80fd5380",
   242 => x"74708405",
   243 => x"560cff13",
   244 => x"53728025",
   245 => x"f238b4f8",
   246 => x"52b39c51",
   247 => x"98bb2d02",
   248 => x"90050d04",
   249 => x"02d8050d",
   250 => x"810bfec4",
   251 => x"0c840bfe",
   252 => x"c40c7b52",
   253 => x"b39c5195",
   254 => x"df2db2fc",
   255 => x"0853b2fc",
   256 => x"08802e81",
   257 => x"c038ae8c",
   258 => x"5185f12d",
   259 => x"b3a00856",
   260 => x"800bff17",
   261 => x"58597679",
   262 => x"2e8b3881",
   263 => x"1977812a",
   264 => x"585976f7",
   265 => x"38f71976",
   266 => x"9fff0654",
   267 => x"5972802e",
   268 => x"8b38fc80",
   269 => x"16b39c52",
   270 => x"5697e82d",
   271 => x"80762580",
   272 => x"fd387852",
   273 => x"76518480",
   274 => x"2db4f852",
   275 => x"b39c5198",
   276 => x"952db2fc",
   277 => x"0853b2fc",
   278 => x"08802e80",
   279 => x"c838b4f8",
   280 => x"5a805889",
   281 => x"92047970",
   282 => x"84055b08",
   283 => x"7083fe80",
   284 => x"0671882b",
   285 => x"83fe8006",
   286 => x"71882a07",
   287 => x"72882a83",
   288 => x"fe800673",
   289 => x"982a07fe",
   290 => x"c80cfec8",
   291 => x"0c568419",
   292 => x"59537553",
   293 => x"84807625",
   294 => x"84388480",
   295 => x"53727824",
   296 => x"c53889ae",
   297 => x"04ae9c51",
   298 => x"85f12d89",
   299 => x"c504b39c",
   300 => x"5197e82d",
   301 => x"fc801681",
   302 => x"18585688",
   303 => x"bc04820b",
   304 => x"fec40c81",
   305 => x"5372b2fc",
   306 => x"0c02a805",
   307 => x"0d04a5a4",
   308 => x"2d0402ec",
   309 => x"050d8117",
   310 => x"54805573",
   311 => x"752ea338",
   312 => x"7451958a",
   313 => x"2db2fc08",
   314 => x"b2fc0809",
   315 => x"810570b2",
   316 => x"fc08079f",
   317 => x"2a767131",
   318 => x"81195957",
   319 => x"51535373",
   320 => x"df387280",
   321 => x"2e983880",
   322 => x"0b8b1481",
   323 => x"b72daeac",
   324 => x"5185f12d",
   325 => x"725185f1",
   326 => x"2d725187",
   327 => x"e42db088",
   328 => x"51a7822d",
   329 => x"a5a42d80",
   330 => x"5184e52d",
   331 => x"0294050d",
   332 => x"0402e805",
   333 => x"0d807056",
   334 => x"5675b2ac",
   335 => x"0825af38",
   336 => x"b9840876",
   337 => x"2ea83874",
   338 => x"51958a2d",
   339 => x"b2fc0809",
   340 => x"810570b2",
   341 => x"fc08079f",
   342 => x"2a770581",
   343 => x"17575752",
   344 => x"75b2ac08",
   345 => x"258838b9",
   346 => x"84087526",
   347 => x"da388056",
   348 => x"74b98408",
   349 => x"2780d038",
   350 => x"7451958a",
   351 => x"2d75842b",
   352 => x"52b2fc08",
   353 => x"802eae38",
   354 => x"b3a81281",
   355 => x"17b2fc08",
   356 => x"5657528a",
   357 => x"53737081",
   358 => x"055580f5",
   359 => x"2d727081",
   360 => x"055481b7",
   361 => x"2dff1353",
   362 => x"728025e9",
   363 => x"38807281",
   364 => x"b72d8bbe",
   365 => x"04b2fc08",
   366 => x"b3a81381",
   367 => x"b72d8115",
   368 => x"558b7625",
   369 => x"ffaa3802",
   370 => x"98050d04",
   371 => x"02fc050d",
   372 => x"725170fd",
   373 => x"2ead3870",
   374 => x"fd248a38",
   375 => x"70fc2e80",
   376 => x"c4388cad",
   377 => x"0470fe2e",
   378 => x"b13870ff",
   379 => x"2e098106",
   380 => x"bc38b2ac",
   381 => x"08517080",
   382 => x"2eb338ff",
   383 => x"11b2ac0c",
   384 => x"8cad04b2",
   385 => x"ac08f005",
   386 => x"70b2ac0c",
   387 => x"51708025",
   388 => x"9c38800b",
   389 => x"b2ac0c8c",
   390 => x"ad04b2ac",
   391 => x"088105b2",
   392 => x"ac0c8cad",
   393 => x"04b2ac08",
   394 => x"9005b2ac",
   395 => x"0c8ab12d",
   396 => x"a5e72d02",
   397 => x"84050d04",
   398 => x"02fc050d",
   399 => x"800bb2ac",
   400 => x"0c8ab12d",
   401 => x"b0f851a7",
   402 => x"822d0284",
   403 => x"050d0402",
   404 => x"f4050d80",
   405 => x"5186922d",
   406 => x"810bfec4",
   407 => x"0c800bfe",
   408 => x"c00c840b",
   409 => x"fec40c83",
   410 => x"0bfecc0c",
   411 => x"a2f22da5",
   412 => x"852da2d7",
   413 => x"2da2d72d",
   414 => x"81f72d81",
   415 => x"5184e52d",
   416 => x"a2d72da2",
   417 => x"d72d8151",
   418 => x"84e52dae",
   419 => x"b85185f1",
   420 => x"2d84529c",
   421 => x"ee2d8ef8",
   422 => x"2db2fc08",
   423 => x"802e8638",
   424 => x"fe528dad",
   425 => x"04ff1252",
   426 => x"718024e7",
   427 => x"3871802e",
   428 => x"80f83886",
   429 => x"c22daed0",
   430 => x"5187e42d",
   431 => x"b2fc0880",
   432 => x"2e8f38b0",
   433 => x"8851a782",
   434 => x"2d805184",
   435 => x"e52d8ddb",
   436 => x"04b2fc08",
   437 => x"518cb82d",
   438 => x"a5912da3",
   439 => x"8a2da792",
   440 => x"2db2fc08",
   441 => x"5386ef2d",
   442 => x"b2fc08fe",
   443 => x"c00c86ef",
   444 => x"2db2fc08",
   445 => x"b398082e",
   446 => x"9c38b2fc",
   447 => x"08b3980c",
   448 => x"84527251",
   449 => x"84e52da2",
   450 => x"d72da2d7",
   451 => x"2dff1252",
   452 => x"718025ee",
   453 => x"3872802e",
   454 => x"89388a0b",
   455 => x"fec40c8d",
   456 => x"db04820b",
   457 => x"fec40c8d",
   458 => x"db04aedc",
   459 => x"5185f12d",
   460 => x"800bb2fc",
   461 => x"0c028c05",
   462 => x"0d0402e8",
   463 => x"050d7779",
   464 => x"7b585555",
   465 => x"80537276",
   466 => x"25a33874",
   467 => x"70810556",
   468 => x"80f52d74",
   469 => x"70810556",
   470 => x"80f52d52",
   471 => x"5271712e",
   472 => x"86388151",
   473 => x"8eef0481",
   474 => x"13538ec6",
   475 => x"04805170",
   476 => x"b2fc0c02",
   477 => x"98050d04",
   478 => x"02d8050d",
   479 => x"800bb980",
   480 => x"0cb4f852",
   481 => x"80519fd6",
   482 => x"2db2fc08",
   483 => x"54b2fc08",
   484 => x"8c38aef0",
   485 => x"5185f12d",
   486 => x"73559493",
   487 => x"04805681",
   488 => x"0bb9a40c",
   489 => x"8853aefc",
   490 => x"52b5ae51",
   491 => x"8eba2db2",
   492 => x"fc08762e",
   493 => x"09810687",
   494 => x"38b2fc08",
   495 => x"b9a40c88",
   496 => x"53af8852",
   497 => x"b5ca518e",
   498 => x"ba2db2fc",
   499 => x"088738b2",
   500 => x"fc08b9a4",
   501 => x"0cb9a408",
   502 => x"802e80f6",
   503 => x"38b8be0b",
   504 => x"80f52db8",
   505 => x"bf0b80f5",
   506 => x"2d71982b",
   507 => x"71902b07",
   508 => x"b8c00b80",
   509 => x"f52d7088",
   510 => x"2b7207b8",
   511 => x"c10b80f5",
   512 => x"2d7107b8",
   513 => x"f60b80f5",
   514 => x"2db8f70b",
   515 => x"80f52d71",
   516 => x"882b0753",
   517 => x"5f54525a",
   518 => x"56575573",
   519 => x"81abaa2e",
   520 => x"0981068d",
   521 => x"387551a0",
   522 => x"f12db2fc",
   523 => x"085690be",
   524 => x"047382d4",
   525 => x"d52e8738",
   526 => x"af945190",
   527 => x"ff04b4f8",
   528 => x"5275519f",
   529 => x"d62db2fc",
   530 => x"0855b2fc",
   531 => x"08802e83",
   532 => x"c2388853",
   533 => x"af8852b5",
   534 => x"ca518eba",
   535 => x"2db2fc08",
   536 => x"8938810b",
   537 => x"b9800c91",
   538 => x"85048853",
   539 => x"aefc52b5",
   540 => x"ae518eba",
   541 => x"2db2fc08",
   542 => x"802e8a38",
   543 => x"afa85185",
   544 => x"f12d91df",
   545 => x"04b8f60b",
   546 => x"80f52d54",
   547 => x"7380d52e",
   548 => x"09810680",
   549 => x"ca38b8f7",
   550 => x"0b80f52d",
   551 => x"547381aa",
   552 => x"2e098106",
   553 => x"ba38800b",
   554 => x"b4f80b80",
   555 => x"f52d5654",
   556 => x"7481e92e",
   557 => x"83388154",
   558 => x"7481eb2e",
   559 => x"8c388055",
   560 => x"73752e09",
   561 => x"810682cb",
   562 => x"38b5830b",
   563 => x"80f52d55",
   564 => x"748d38b5",
   565 => x"840b80f5",
   566 => x"2d547382",
   567 => x"2e863880",
   568 => x"55949304",
   569 => x"b5850b80",
   570 => x"f52d70b8",
   571 => x"f80cff05",
   572 => x"b8fc0cb5",
   573 => x"860b80f5",
   574 => x"2db5870b",
   575 => x"80f52d58",
   576 => x"76057782",
   577 => x"80290570",
   578 => x"b9880cb5",
   579 => x"880b80f5",
   580 => x"2d70b99c",
   581 => x"0cb98008",
   582 => x"59575876",
   583 => x"802e81a3",
   584 => x"388853af",
   585 => x"8852b5ca",
   586 => x"518eba2d",
   587 => x"b2fc0881",
   588 => x"e238b8f8",
   589 => x"0870842b",
   590 => x"b9840c70",
   591 => x"b9980cb5",
   592 => x"9d0b80f5",
   593 => x"2db59c0b",
   594 => x"80f52d71",
   595 => x"82802905",
   596 => x"b59e0b80",
   597 => x"f52d7084",
   598 => x"80802912",
   599 => x"b59f0b80",
   600 => x"f52d7081",
   601 => x"800a2912",
   602 => x"70b9a00c",
   603 => x"b99c0871",
   604 => x"29b98808",
   605 => x"0570b98c",
   606 => x"0cb5a50b",
   607 => x"80f52db5",
   608 => x"a40b80f5",
   609 => x"2d718280",
   610 => x"2905b5a6",
   611 => x"0b80f52d",
   612 => x"70848080",
   613 => x"2912b5a7",
   614 => x"0b80f52d",
   615 => x"70982b81",
   616 => x"f00a0672",
   617 => x"0570b990",
   618 => x"0cfe117e",
   619 => x"297705b9",
   620 => x"940c5259",
   621 => x"5243545e",
   622 => x"51525952",
   623 => x"5d575957",
   624 => x"949104b5",
   625 => x"8a0b80f5",
   626 => x"2db5890b",
   627 => x"80f52d71",
   628 => x"82802905",
   629 => x"70b9840c",
   630 => x"70a02983",
   631 => x"ff057089",
   632 => x"2a70b998",
   633 => x"0cb58f0b",
   634 => x"80f52db5",
   635 => x"8e0b80f5",
   636 => x"2d718280",
   637 => x"290570b9",
   638 => x"a00c7b71",
   639 => x"291e70b9",
   640 => x"940c7db9",
   641 => x"900c7305",
   642 => x"b98c0c55",
   643 => x"5e515155",
   644 => x"55815574",
   645 => x"b2fc0c02",
   646 => x"a8050d04",
   647 => x"02ec050d",
   648 => x"7670872c",
   649 => x"7180ff06",
   650 => x"555654b9",
   651 => x"80088a38",
   652 => x"73882c74",
   653 => x"81ff0654",
   654 => x"55b4f852",
   655 => x"b9880815",
   656 => x"519fd62d",
   657 => x"b2fc0854",
   658 => x"b2fc0880",
   659 => x"2eb338b9",
   660 => x"8008802e",
   661 => x"98387284",
   662 => x"29b4f805",
   663 => x"70085253",
   664 => x"a0f12db2",
   665 => x"fc08f00a",
   666 => x"065394ff",
   667 => x"047210b4",
   668 => x"f8057080",
   669 => x"e02d5253",
   670 => x"a1a12db2",
   671 => x"fc085372",
   672 => x"5473b2fc",
   673 => x"0c029405",
   674 => x"0d0402ec",
   675 => x"050d7670",
   676 => x"842cb994",
   677 => x"0805718f",
   678 => x"06525553",
   679 => x"728938b4",
   680 => x"f8527351",
   681 => x"9fd62d72",
   682 => x"a029b4f8",
   683 => x"05548074",
   684 => x"80f52d54",
   685 => x"5572752e",
   686 => x"83388155",
   687 => x"7281e52e",
   688 => x"93387480",
   689 => x"2e8e388b",
   690 => x"1480f52d",
   691 => x"98065372",
   692 => x"802e8338",
   693 => x"805473b2",
   694 => x"fc0c0294",
   695 => x"050d0402",
   696 => x"cc050d7e",
   697 => x"605e5a80",
   698 => x"0bb99008",
   699 => x"b9940859",
   700 => x"5c568058",
   701 => x"b9840878",
   702 => x"2e81ae38",
   703 => x"778f06a0",
   704 => x"17575473",
   705 => x"8f38b4f8",
   706 => x"52765181",
   707 => x"17579fd6",
   708 => x"2db4f856",
   709 => x"807680f5",
   710 => x"2d565474",
   711 => x"742e8338",
   712 => x"81547481",
   713 => x"e52e80f6",
   714 => x"38817075",
   715 => x"06555c73",
   716 => x"802e80ea",
   717 => x"388b1680",
   718 => x"f52d9806",
   719 => x"597880de",
   720 => x"388b537c",
   721 => x"5275518e",
   722 => x"ba2db2fc",
   723 => x"0880cf38",
   724 => x"9c160851",
   725 => x"a0f12db2",
   726 => x"fc08841b",
   727 => x"0c9a1680",
   728 => x"e02d51a1",
   729 => x"a12db2fc",
   730 => x"08b2fc08",
   731 => x"881c0cb2",
   732 => x"fc085555",
   733 => x"b9800880",
   734 => x"2e983894",
   735 => x"1680e02d",
   736 => x"51a1a12d",
   737 => x"b2fc0890",
   738 => x"2b83fff0",
   739 => x"0a067016",
   740 => x"51547388",
   741 => x"1b0c787a",
   742 => x"0c7b5497",
   743 => x"df048118",
   744 => x"58b98408",
   745 => x"7826fed4",
   746 => x"38b98008",
   747 => x"802eae38",
   748 => x"7a51949c",
   749 => x"2db2fc08",
   750 => x"b2fc0880",
   751 => x"fffffff8",
   752 => x"06555b73",
   753 => x"80ffffff",
   754 => x"f82e9238",
   755 => x"b2fc08fe",
   756 => x"05b8f808",
   757 => x"29b98c08",
   758 => x"055795f2",
   759 => x"04805473",
   760 => x"b2fc0c02",
   761 => x"b4050d04",
   762 => x"02f4050d",
   763 => x"74700881",
   764 => x"05710c70",
   765 => x"08b8fc08",
   766 => x"06535371",
   767 => x"8e388813",
   768 => x"0851949c",
   769 => x"2db2fc08",
   770 => x"88140c81",
   771 => x"0bb2fc0c",
   772 => x"028c050d",
   773 => x"0402f005",
   774 => x"0d758811",
   775 => x"08fe05b8",
   776 => x"f80829b9",
   777 => x"8c081172",
   778 => x"08b8fc08",
   779 => x"06057955",
   780 => x"5354549f",
   781 => x"d62d0290",
   782 => x"050d0402",
   783 => x"f0050d75",
   784 => x"881108fe",
   785 => x"05b8f808",
   786 => x"29b98c08",
   787 => x"117208b8",
   788 => x"fc080605",
   789 => x"79555354",
   790 => x"549e962d",
   791 => x"0290050d",
   792 => x"0402f405",
   793 => x"0dd45281",
   794 => x"ff720c71",
   795 => x"085381ff",
   796 => x"720c7288",
   797 => x"2b83fe80",
   798 => x"06720870",
   799 => x"81ff0651",
   800 => x"525381ff",
   801 => x"720c7271",
   802 => x"07882b72",
   803 => x"087081ff",
   804 => x"06515253",
   805 => x"81ff720c",
   806 => x"72710788",
   807 => x"2b720870",
   808 => x"81ff0672",
   809 => x"07b2fc0c",
   810 => x"5253028c",
   811 => x"050d0402",
   812 => x"f4050d74",
   813 => x"767181ff",
   814 => x"06d40c53",
   815 => x"53b9a808",
   816 => x"85387189",
   817 => x"2b527198",
   818 => x"2ad40c71",
   819 => x"902a7081",
   820 => x"ff06d40c",
   821 => x"5171882a",
   822 => x"7081ff06",
   823 => x"d40c5171",
   824 => x"81ff06d4",
   825 => x"0c72902a",
   826 => x"7081ff06",
   827 => x"d40c51d4",
   828 => x"087081ff",
   829 => x"06515182",
   830 => x"b8bf5270",
   831 => x"81ff2e09",
   832 => x"81069438",
   833 => x"81ff0bd4",
   834 => x"0cd40870",
   835 => x"81ff06ff",
   836 => x"14545151",
   837 => x"71e53870",
   838 => x"b2fc0c02",
   839 => x"8c050d04",
   840 => x"02fc050d",
   841 => x"81c75181",
   842 => x"ff0bd40c",
   843 => x"ff115170",
   844 => x"8025f438",
   845 => x"0284050d",
   846 => x"0402f005",
   847 => x"0d9aa02d",
   848 => x"8fcf5380",
   849 => x"5287fc80",
   850 => x"f75199af",
   851 => x"2db2fc08",
   852 => x"54b2fc08",
   853 => x"812e0981",
   854 => x"06a33881",
   855 => x"ff0bd40c",
   856 => x"820a5284",
   857 => x"9c80e951",
   858 => x"99af2db2",
   859 => x"fc088b38",
   860 => x"81ff0bd4",
   861 => x"0c73539b",
   862 => x"83049aa0",
   863 => x"2dff1353",
   864 => x"72c13872",
   865 => x"b2fc0c02",
   866 => x"90050d04",
   867 => x"02f4050d",
   868 => x"81ff0bd4",
   869 => x"0c935380",
   870 => x"5287fc80",
   871 => x"c15199af",
   872 => x"2db2fc08",
   873 => x"8b3881ff",
   874 => x"0bd40c81",
   875 => x"539bb904",
   876 => x"9aa02dff",
   877 => x"135372df",
   878 => x"3872b2fc",
   879 => x"0c028c05",
   880 => x"0d0402f0",
   881 => x"050d9aa0",
   882 => x"2d83aa52",
   883 => x"849c80c8",
   884 => x"5199af2d",
   885 => x"b2fc0881",
   886 => x"2e098106",
   887 => x"923898e1",
   888 => x"2db2fc08",
   889 => x"83ffff06",
   890 => x"537283aa",
   891 => x"2e97389b",
   892 => x"8c2d9c80",
   893 => x"0481549c",
   894 => x"e504afb4",
   895 => x"5185f12d",
   896 => x"80549ce5",
   897 => x"0481ff0b",
   898 => x"d40cb153",
   899 => x"9ab92db2",
   900 => x"fc08802e",
   901 => x"80c03880",
   902 => x"5287fc80",
   903 => x"fa5199af",
   904 => x"2db2fc08",
   905 => x"b13881ff",
   906 => x"0bd40cd4",
   907 => x"085381ff",
   908 => x"0bd40c81",
   909 => x"ff0bd40c",
   910 => x"81ff0bd4",
   911 => x"0c81ff0b",
   912 => x"d40c7286",
   913 => x"2a708106",
   914 => x"b2fc0856",
   915 => x"51537280",
   916 => x"2e93389b",
   917 => x"f5047282",
   918 => x"2eff9f38",
   919 => x"ff135372",
   920 => x"ffaa3872",
   921 => x"5473b2fc",
   922 => x"0c029005",
   923 => x"0d0402f0",
   924 => x"050d810b",
   925 => x"b9a80c84",
   926 => x"54d00870",
   927 => x"8f2a7081",
   928 => x"06515153",
   929 => x"72f33872",
   930 => x"d00c9aa0",
   931 => x"2dafc451",
   932 => x"85f12dd0",
   933 => x"08708f2a",
   934 => x"70810651",
   935 => x"515372f3",
   936 => x"38810bd0",
   937 => x"0cb15380",
   938 => x"5284d480",
   939 => x"c05199af",
   940 => x"2db2fc08",
   941 => x"812ea138",
   942 => x"72822e09",
   943 => x"81068c38",
   944 => x"afd05185",
   945 => x"f12d8053",
   946 => x"9e8d04ff",
   947 => x"135372d7",
   948 => x"38ff1454",
   949 => x"73ffa238",
   950 => x"9bc22db2",
   951 => x"fc08b9a8",
   952 => x"0cb2fc08",
   953 => x"8b388152",
   954 => x"87fc80d0",
   955 => x"5199af2d",
   956 => x"81ff0bd4",
   957 => x"0cd00870",
   958 => x"8f2a7081",
   959 => x"06515153",
   960 => x"72f33872",
   961 => x"d00c81ff",
   962 => x"0bd40c81",
   963 => x"5372b2fc",
   964 => x"0c029005",
   965 => x"0d0402e8",
   966 => x"050d7856",
   967 => x"81ff0bd4",
   968 => x"0cd00870",
   969 => x"8f2a7081",
   970 => x"06515153",
   971 => x"72f33882",
   972 => x"810bd00c",
   973 => x"81ff0bd4",
   974 => x"0c775287",
   975 => x"fc80d851",
   976 => x"99af2db2",
   977 => x"fc08802e",
   978 => x"8c38afe8",
   979 => x"5185f12d",
   980 => x"81539fcd",
   981 => x"0481ff0b",
   982 => x"d40c81fe",
   983 => x"0bd40c80",
   984 => x"ff557570",
   985 => x"84055708",
   986 => x"70982ad4",
   987 => x"0c70902c",
   988 => x"7081ff06",
   989 => x"d40c5470",
   990 => x"882c7081",
   991 => x"ff06d40c",
   992 => x"547081ff",
   993 => x"06d40c54",
   994 => x"ff155574",
   995 => x"8025d338",
   996 => x"81ff0bd4",
   997 => x"0c81ff0b",
   998 => x"d40c81ff",
   999 => x"0bd40c86",
  1000 => x"8da05481",
  1001 => x"ff0bd40c",
  1002 => x"d40881ff",
  1003 => x"06557487",
  1004 => x"38ff1454",
  1005 => x"73ed3881",
  1006 => x"ff0bd40c",
  1007 => x"d008708f",
  1008 => x"2a708106",
  1009 => x"51515372",
  1010 => x"f33872d0",
  1011 => x"0c72b2fc",
  1012 => x"0c029805",
  1013 => x"0d0402e8",
  1014 => x"050d7855",
  1015 => x"805681ff",
  1016 => x"0bd40cd0",
  1017 => x"08708f2a",
  1018 => x"70810651",
  1019 => x"515372f3",
  1020 => x"3882810b",
  1021 => x"d00c81ff",
  1022 => x"0bd40c77",
  1023 => x"5287fc80",
  1024 => x"d15199af",
  1025 => x"2d80dbc6",
  1026 => x"df54b2fc",
  1027 => x"08802e8a",
  1028 => x"38ae9c51",
  1029 => x"85f12da0",
  1030 => x"e80481ff",
  1031 => x"0bd40cd4",
  1032 => x"087081ff",
  1033 => x"06515372",
  1034 => x"81fe2e09",
  1035 => x"81069d38",
  1036 => x"80ff5398",
  1037 => x"e12db2fc",
  1038 => x"08757084",
  1039 => x"05570cff",
  1040 => x"13537280",
  1041 => x"25ed3881",
  1042 => x"56a0d204",
  1043 => x"ff145473",
  1044 => x"c93881ff",
  1045 => x"0bd40cd0",
  1046 => x"08708f2a",
  1047 => x"70810651",
  1048 => x"515372f3",
  1049 => x"3872d00c",
  1050 => x"75b2fc0c",
  1051 => x"0298050d",
  1052 => x"0402f405",
  1053 => x"0d747088",
  1054 => x"2a83fe80",
  1055 => x"06707298",
  1056 => x"2a077288",
  1057 => x"2b87fc80",
  1058 => x"80067398",
  1059 => x"2b81f00a",
  1060 => x"06717307",
  1061 => x"07b2fc0c",
  1062 => x"56515351",
  1063 => x"028c050d",
  1064 => x"0402f805",
  1065 => x"0d028e05",
  1066 => x"80f52d74",
  1067 => x"882b0770",
  1068 => x"83ffff06",
  1069 => x"b2fc0c51",
  1070 => x"0288050d",
  1071 => x"0402fc05",
  1072 => x"0d725180",
  1073 => x"710c800b",
  1074 => x"84120c02",
  1075 => x"84050d04",
  1076 => x"02f0050d",
  1077 => x"75700884",
  1078 => x"12085353",
  1079 => x"53ff5471",
  1080 => x"712ea838",
  1081 => x"a58b2d84",
  1082 => x"13087084",
  1083 => x"29148811",
  1084 => x"70087081",
  1085 => x"ff068418",
  1086 => x"08811187",
  1087 => x"06841a0c",
  1088 => x"53515551",
  1089 => x"5151a585",
  1090 => x"2d715473",
  1091 => x"b2fc0c02",
  1092 => x"90050d04",
  1093 => x"02f8050d",
  1094 => x"a58b2de0",
  1095 => x"08708b2a",
  1096 => x"70810651",
  1097 => x"52527080",
  1098 => x"2e9d38b9",
  1099 => x"ac087084",
  1100 => x"29b9b405",
  1101 => x"7381ff06",
  1102 => x"710c5151",
  1103 => x"b9ac0881",
  1104 => x"118706b9",
  1105 => x"ac0c5180",
  1106 => x"0bb9d40c",
  1107 => x"a4fe2da5",
  1108 => x"852d0288",
  1109 => x"050d0402",
  1110 => x"fc050da5",
  1111 => x"8b2d810b",
  1112 => x"b9d40ca5",
  1113 => x"852db9d4",
  1114 => x"085170fa",
  1115 => x"38028405",
  1116 => x"0d0402fc",
  1117 => x"050db9ac",
  1118 => x"51a1bd2d",
  1119 => x"a29451a4",
  1120 => x"fa2da4a4",
  1121 => x"2d028405",
  1122 => x"0d0402f4",
  1123 => x"050da48c",
  1124 => x"04b2fc08",
  1125 => x"81f02e09",
  1126 => x"81068938",
  1127 => x"810bb2f0",
  1128 => x"0ca48c04",
  1129 => x"b2fc0881",
  1130 => x"e02e0981",
  1131 => x"06893881",
  1132 => x"0bb2f40c",
  1133 => x"a48c04b2",
  1134 => x"fc0852b2",
  1135 => x"f408802e",
  1136 => x"8838b2fc",
  1137 => x"08818005",
  1138 => x"5271842c",
  1139 => x"728f0653",
  1140 => x"53b2f008",
  1141 => x"802e9938",
  1142 => x"728429b2",
  1143 => x"b0057213",
  1144 => x"81712b70",
  1145 => x"09730806",
  1146 => x"730c5153",
  1147 => x"53a48204",
  1148 => x"728429b2",
  1149 => x"b0057213",
  1150 => x"83712b72",
  1151 => x"0807720c",
  1152 => x"5353800b",
  1153 => x"b2f40c80",
  1154 => x"0bb2f00c",
  1155 => x"b9ac51a1",
  1156 => x"d02db2fc",
  1157 => x"08ff24fe",
  1158 => x"f838800b",
  1159 => x"b2fc0c02",
  1160 => x"8c050d04",
  1161 => x"02f8050d",
  1162 => x"b2b0528f",
  1163 => x"51807270",
  1164 => x"8405540c",
  1165 => x"ff115170",
  1166 => x"8025f238",
  1167 => x"0288050d",
  1168 => x"0402f005",
  1169 => x"0d7551a5",
  1170 => x"8b2d7082",
  1171 => x"2cfc06b2",
  1172 => x"b0117210",
  1173 => x"9e067108",
  1174 => x"70722a70",
  1175 => x"83068274",
  1176 => x"2b700974",
  1177 => x"06760c54",
  1178 => x"51565753",
  1179 => x"5153a585",
  1180 => x"2d71b2fc",
  1181 => x"0c029005",
  1182 => x"0d047198",
  1183 => x"0c04ffb0",
  1184 => x"08b2fc0c",
  1185 => x"04810bff",
  1186 => x"b00c0480",
  1187 => x"0bffb00c",
  1188 => x"0402fc05",
  1189 => x"0d810bb2",
  1190 => x"f80c8151",
  1191 => x"84e52d02",
  1192 => x"84050d04",
  1193 => x"02fc050d",
  1194 => x"800bb2f8",
  1195 => x"0c805184",
  1196 => x"e52d0284",
  1197 => x"050d0402",
  1198 => x"ec050d76",
  1199 => x"54805287",
  1200 => x"0b881580",
  1201 => x"f52d5653",
  1202 => x"74722483",
  1203 => x"38a05372",
  1204 => x"5182ee2d",
  1205 => x"81128b15",
  1206 => x"80f52d54",
  1207 => x"52727225",
  1208 => x"de380294",
  1209 => x"050d0402",
  1210 => x"f0050db9",
  1211 => x"dc085481",
  1212 => x"f72d800b",
  1213 => x"b9e00c73",
  1214 => x"08802e81",
  1215 => x"8038820b",
  1216 => x"b3900cb9",
  1217 => x"e0088f06",
  1218 => x"b38c0c73",
  1219 => x"08527183",
  1220 => x"2e963871",
  1221 => x"83268938",
  1222 => x"71812eaf",
  1223 => x"38a6e804",
  1224 => x"71852e9f",
  1225 => x"38a6e804",
  1226 => x"881480f5",
  1227 => x"2d841508",
  1228 => x"aff85354",
  1229 => x"5285f12d",
  1230 => x"71842913",
  1231 => x"70085252",
  1232 => x"a6ec0473",
  1233 => x"51a5b72d",
  1234 => x"a6e804b9",
  1235 => x"d8088815",
  1236 => x"082c7081",
  1237 => x"06515271",
  1238 => x"802e8738",
  1239 => x"affc51a6",
  1240 => x"e504b080",
  1241 => x"5185f12d",
  1242 => x"84140851",
  1243 => x"85f12db9",
  1244 => x"e0088105",
  1245 => x"b9e00c8c",
  1246 => x"1454a5f7",
  1247 => x"04029005",
  1248 => x"0d0471b9",
  1249 => x"dc0ca5e7",
  1250 => x"2db9e008",
  1251 => x"ff05b9e4",
  1252 => x"0c0402ec",
  1253 => x"050db9dc",
  1254 => x"085580f8",
  1255 => x"51a4c12d",
  1256 => x"b2fc0881",
  1257 => x"2a708106",
  1258 => x"5152719b",
  1259 => x"388751a4",
  1260 => x"c12db2fc",
  1261 => x"08812a70",
  1262 => x"81065152",
  1263 => x"71802eb1",
  1264 => x"38a7c704",
  1265 => x"a38a2d87",
  1266 => x"51a4c12d",
  1267 => x"b2fc08f4",
  1268 => x"38a7d704",
  1269 => x"a38a2d80",
  1270 => x"f851a4c1",
  1271 => x"2db2fc08",
  1272 => x"f338b2f8",
  1273 => x"08813270",
  1274 => x"b2f80c70",
  1275 => x"525284e5",
  1276 => x"2db2f808",
  1277 => x"ae3880da",
  1278 => x"51a4c12d",
  1279 => x"81f551a4",
  1280 => x"c12d81f2",
  1281 => x"51a4c12d",
  1282 => x"81eb51a4",
  1283 => x"c12d81f4",
  1284 => x"51a4c12d",
  1285 => x"81fd51a4",
  1286 => x"c12d81fa",
  1287 => x"51a4c12d",
  1288 => x"acde0481",
  1289 => x"f551a4c1",
  1290 => x"2db2fc08",
  1291 => x"812a7081",
  1292 => x"06515271",
  1293 => x"802eaf38",
  1294 => x"b9e40852",
  1295 => x"71802e89",
  1296 => x"38ff12b9",
  1297 => x"e40ca8e6",
  1298 => x"04b9e008",
  1299 => x"10b9e008",
  1300 => x"05708429",
  1301 => x"16515288",
  1302 => x"1208802e",
  1303 => x"8938ff51",
  1304 => x"88120852",
  1305 => x"712d81f2",
  1306 => x"51a4c12d",
  1307 => x"b2fc0881",
  1308 => x"2a708106",
  1309 => x"51527180",
  1310 => x"2eb138b9",
  1311 => x"e008ff11",
  1312 => x"b9e40856",
  1313 => x"53537372",
  1314 => x"25893881",
  1315 => x"14b9e40c",
  1316 => x"a9ab0472",
  1317 => x"10137084",
  1318 => x"29165152",
  1319 => x"88120880",
  1320 => x"2e8938fe",
  1321 => x"51881208",
  1322 => x"52712d81",
  1323 => x"fd51a4c1",
  1324 => x"2db2fc08",
  1325 => x"812a7081",
  1326 => x"06515271",
  1327 => x"802e8638",
  1328 => x"800bb9e4",
  1329 => x"0c81fa51",
  1330 => x"a4c12db2",
  1331 => x"fc08812a",
  1332 => x"70810651",
  1333 => x"5271802e",
  1334 => x"8938b9e0",
  1335 => x"08ff05b9",
  1336 => x"e40cb9e4",
  1337 => x"08705354",
  1338 => x"73802e8a",
  1339 => x"388c15ff",
  1340 => x"155555a9",
  1341 => x"e804820b",
  1342 => x"b3900c71",
  1343 => x"8f06b38c",
  1344 => x"0c81eb51",
  1345 => x"a4c12db2",
  1346 => x"fc08812a",
  1347 => x"70810651",
  1348 => x"5271802e",
  1349 => x"ad387408",
  1350 => x"852e0981",
  1351 => x"06a43888",
  1352 => x"1580f52d",
  1353 => x"ff055271",
  1354 => x"881681b7",
  1355 => x"2d71982b",
  1356 => x"52718025",
  1357 => x"8838800b",
  1358 => x"881681b7",
  1359 => x"2d7451a5",
  1360 => x"b72d81f4",
  1361 => x"51a4c12d",
  1362 => x"b2fc0881",
  1363 => x"2a708106",
  1364 => x"51527180",
  1365 => x"2eb33874",
  1366 => x"08852e09",
  1367 => x"8106aa38",
  1368 => x"881580f5",
  1369 => x"2d810552",
  1370 => x"71881681",
  1371 => x"b72d7181",
  1372 => x"ff068b16",
  1373 => x"80f52d54",
  1374 => x"52727227",
  1375 => x"87387288",
  1376 => x"1681b72d",
  1377 => x"7451a5b7",
  1378 => x"2d80da51",
  1379 => x"a4c12db2",
  1380 => x"fc08812a",
  1381 => x"70810651",
  1382 => x"5271802e",
  1383 => x"80ff38b9",
  1384 => x"dc08b9e4",
  1385 => x"08555373",
  1386 => x"802e8a38",
  1387 => x"8c13ff15",
  1388 => x"5553aba7",
  1389 => x"04720852",
  1390 => x"71822ea6",
  1391 => x"38718226",
  1392 => x"89387181",
  1393 => x"2ea938ac",
  1394 => x"9d047183",
  1395 => x"2eb13871",
  1396 => x"842e0981",
  1397 => x"0680c638",
  1398 => x"88130851",
  1399 => x"a7822dac",
  1400 => x"9d04b9e4",
  1401 => x"08518813",
  1402 => x"0852712d",
  1403 => x"ac9d0481",
  1404 => x"0b881408",
  1405 => x"2bb9d808",
  1406 => x"32b9d80c",
  1407 => x"ac9a0488",
  1408 => x"1380f52d",
  1409 => x"81058b14",
  1410 => x"80f52d53",
  1411 => x"54717424",
  1412 => x"83388054",
  1413 => x"73881481",
  1414 => x"b72da5e7",
  1415 => x"2d805480",
  1416 => x"0bb3900c",
  1417 => x"738f06b3",
  1418 => x"8c0ca052",
  1419 => x"73b9e408",
  1420 => x"2e098106",
  1421 => x"9838b9e0",
  1422 => x"08ff0574",
  1423 => x"32700981",
  1424 => x"05707207",
  1425 => x"9f2a9171",
  1426 => x"31515153",
  1427 => x"53715182",
  1428 => x"ee2d8114",
  1429 => x"548e7425",
  1430 => x"c638b2f8",
  1431 => x"085271b2",
  1432 => x"fc0c0294",
  1433 => x"050d0400",
  1434 => x"00ffffff",
  1435 => x"ff00ffff",
  1436 => x"ffff00ff",
  1437 => x"ffffff00",
  1438 => x"52657365",
  1439 => x"74000000",
  1440 => x"53617665",
  1441 => x"20736574",
  1442 => x"74696e67",
  1443 => x"73000000",
  1444 => x"5363616e",
  1445 => x"6c696e65",
  1446 => x"73000000",
  1447 => x"4c6f6164",
  1448 => x"20524f4d",
  1449 => x"20100000",
  1450 => x"45786974",
  1451 => x"00000000",
  1452 => x"50432045",
  1453 => x"6e67696e",
  1454 => x"65206d6f",
  1455 => x"64650000",
  1456 => x"54757262",
  1457 => x"6f677261",
  1458 => x"66782031",
  1459 => x"36206d6f",
  1460 => x"64650000",
  1461 => x"56474120",
  1462 => x"2d203331",
  1463 => x"4b487a2c",
  1464 => x"20363048",
  1465 => x"7a000000",
  1466 => x"5456202d",
  1467 => x"20343830",
  1468 => x"692c2036",
  1469 => x"30487a00",
  1470 => x"4261636b",
  1471 => x"00000000",
  1472 => x"46504741",
  1473 => x"50434520",
  1474 => x"43464700",
  1475 => x"4c6f6164",
  1476 => x"696e6720",
  1477 => x"524f4d0a",
  1478 => x"00000000",
  1479 => x"52656164",
  1480 => x"20666169",
  1481 => x"6c65640a",
  1482 => x"00000000",
  1483 => x"4c6f6164",
  1484 => x"696e6720",
  1485 => x"00000000",
  1486 => x"496e6974",
  1487 => x"69616c69",
  1488 => x"7a696e67",
  1489 => x"20534420",
  1490 => x"63617264",
  1491 => x"0a000000",
  1492 => x"424f4f54",
  1493 => x"20202020",
  1494 => x"50434500",
  1495 => x"43617264",
  1496 => x"20696e69",
  1497 => x"74206661",
  1498 => x"696c6564",
  1499 => x"0a000000",
  1500 => x"4d425220",
  1501 => x"6661696c",
  1502 => x"0a000000",
  1503 => x"46415431",
  1504 => x"36202020",
  1505 => x"00000000",
  1506 => x"46415433",
  1507 => x"32202020",
  1508 => x"00000000",
  1509 => x"4e6f2070",
  1510 => x"61727469",
  1511 => x"74696f6e",
  1512 => x"20736967",
  1513 => x"0a000000",
  1514 => x"42616420",
  1515 => x"70617274",
  1516 => x"0a000000",
  1517 => x"53444843",
  1518 => x"20657272",
  1519 => x"6f72210a",
  1520 => x"00000000",
  1521 => x"53442069",
  1522 => x"6e69742e",
  1523 => x"2e2e0a00",
  1524 => x"53442063",
  1525 => x"61726420",
  1526 => x"72657365",
  1527 => x"74206661",
  1528 => x"696c6564",
  1529 => x"210a0000",
  1530 => x"57726974",
  1531 => x"65206661",
  1532 => x"696c6564",
  1533 => x"0a000000",
  1534 => x"16200000",
  1535 => x"14200000",
  1536 => x"15200000",
  1537 => x"00000002",
  1538 => x"00000002",
  1539 => x"00001678",
  1540 => x"000004ce",
  1541 => x"00000002",
  1542 => x"00001680",
  1543 => x"000003a2",
  1544 => x"00000003",
  1545 => x"00001870",
  1546 => x"00000002",
  1547 => x"00000001",
  1548 => x"00001690",
  1549 => x"00000001",
  1550 => x"00000003",
  1551 => x"00001868",
  1552 => x"00000002",
  1553 => x"00000002",
  1554 => x"0000169c",
  1555 => x"00000638",
  1556 => x"00000002",
  1557 => x"000016a8",
  1558 => x"000012a4",
  1559 => x"00000000",
  1560 => x"00000000",
  1561 => x"00000000",
  1562 => x"000016b0",
  1563 => x"000016c0",
  1564 => x"000016d4",
  1565 => x"000016e8",
  1566 => x"00000002",
  1567 => x"000019a8",
  1568 => x"000004d2",
  1569 => x"00000002",
  1570 => x"000019b8",
  1571 => x"000004d2",
  1572 => x"00000002",
  1573 => x"000019c8",
  1574 => x"000004d2",
  1575 => x"00000002",
  1576 => x"000019d8",
  1577 => x"000004d2",
  1578 => x"00000002",
  1579 => x"000019e8",
  1580 => x"000004d2",
  1581 => x"00000002",
  1582 => x"000019f8",
  1583 => x"000004d2",
  1584 => x"00000002",
  1585 => x"00001a08",
  1586 => x"000004d2",
  1587 => x"00000002",
  1588 => x"00001a18",
  1589 => x"000004d2",
  1590 => x"00000002",
  1591 => x"00001a28",
  1592 => x"000004d2",
  1593 => x"00000002",
  1594 => x"00001a38",
  1595 => x"000004d2",
  1596 => x"00000002",
  1597 => x"00001a48",
  1598 => x"000004d2",
  1599 => x"00000002",
  1600 => x"00001a58",
  1601 => x"000004d2",
  1602 => x"00000002",
  1603 => x"00001a68",
  1604 => x"000004d2",
  1605 => x"00000004",
  1606 => x"000016f8",
  1607 => x"00001808",
  1608 => x"00000000",
  1609 => x"00000000",
  1610 => x"000005cc",
  1611 => x"00000000",
  1612 => x"00000000",
  1613 => x"00000000",
  1614 => x"00000000",
  1615 => x"00000000",
  1616 => x"00000000",
  1617 => x"00000000",
  1618 => x"00000000",
  1619 => x"00000000",
  1620 => x"00000000",
  1621 => x"00000000",
  1622 => x"00000000",
  1623 => x"00000000",
  1624 => x"00000000",
  1625 => x"00000000",
  1626 => x"00000000",
  1627 => x"00000000",
  1628 => x"00000000",
  1629 => x"00000000",
  1630 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

