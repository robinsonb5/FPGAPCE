-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb6",
     9 => x"b0080b0b",
    10 => x"0bb6b408",
    11 => x"0b0b0bb6",
    12 => x"b8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b6b80c0b",
    16 => x"0b0bb6b4",
    17 => x"0c0b0b0b",
    18 => x"b6b00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb0a0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b6b070bd",
    57 => x"ac278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"8d860402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b6c00c9f",
    65 => x"0bb6c40c",
    66 => x"a0717081",
    67 => x"055334b6",
    68 => x"c408ff05",
    69 => x"b6c40cb6",
    70 => x"c4088025",
    71 => x"eb38b6c0",
    72 => x"08ff05b6",
    73 => x"c00cb6c0",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0bb6c0",
    94 => x"08258f38",
    95 => x"82b22db6",
    96 => x"c008ff05",
    97 => x"b6c00c82",
    98 => x"f404b6c0",
    99 => x"08b6c408",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38b6c008",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134b6",
   108 => x"c4088105",
   109 => x"b6c40cb6",
   110 => x"c408519f",
   111 => x"7125e238",
   112 => x"800bb6c4",
   113 => x"0cb6c008",
   114 => x"8105b6c0",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"b6c40881",
   120 => x"05b6c40c",
   121 => x"b6c408a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"b6c40cb6",
   125 => x"c0088105",
   126 => x"b6c00c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800bb6",
   155 => x"c80cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820bb6c8",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"b6c80884",
   167 => x"07b6c80c",
   168 => x"5573842b",
   169 => x"87e87125",
   170 => x"83713170",
   171 => x"0b0b0bb3",
   172 => x"a00c8171",
   173 => x"2bf6880c",
   174 => x"fea413ff",
   175 => x"122c7888",
   176 => x"29ff9405",
   177 => x"70812cb6",
   178 => x"c8085258",
   179 => x"52555152",
   180 => x"5476802e",
   181 => x"85387081",
   182 => x"075170f6",
   183 => x"940c7109",
   184 => x"8105f680",
   185 => x"0c720981",
   186 => x"05f6840c",
   187 => x"0294050d",
   188 => x"0402f405",
   189 => x"0d745372",
   190 => x"70810554",
   191 => x"80f52d52",
   192 => x"71802e89",
   193 => x"38715182",
   194 => x"ee2d85f7",
   195 => x"04028c05",
   196 => x"0d0402f4",
   197 => x"050d7470",
   198 => x"8206bd90",
   199 => x"0cb3bc71",
   200 => x"81065454",
   201 => x"51718814",
   202 => x"81b72d70",
   203 => x"822a7081",
   204 => x"06515170",
   205 => x"a01481b7",
   206 => x"2d70b6b0",
   207 => x"0c028c05",
   208 => x"0d0402f8",
   209 => x"050db1b8",
   210 => x"52b6cc51",
   211 => x"96a42db6",
   212 => x"b008802e",
   213 => x"9d38b8b0",
   214 => x"52b6cc51",
   215 => x"98da2db8",
   216 => x"b008b6d8",
   217 => x"0cb8b008",
   218 => x"fec00cb8",
   219 => x"b0085186",
   220 => x"922d0288",
   221 => x"050d0402",
   222 => x"f0050db1",
   223 => x"b852b6cc",
   224 => x"5196a42d",
   225 => x"b6b00880",
   226 => x"2ea538b6",
   227 => x"d808b8b0",
   228 => x"0cb8b454",
   229 => x"80fd5380",
   230 => x"74708405",
   231 => x"560cff13",
   232 => x"53728025",
   233 => x"f238b8b0",
   234 => x"52b6cc51",
   235 => x"99802d02",
   236 => x"90050d04",
   237 => x"02d4050d",
   238 => x"810bfec4",
   239 => x"0c840bfe",
   240 => x"c40c7c52",
   241 => x"b6cc5196",
   242 => x"a42db6b0",
   243 => x"0853b6b0",
   244 => x"08802e81",
   245 => x"cc38b6d0",
   246 => x"0856800b",
   247 => x"ff175859",
   248 => x"76792e8b",
   249 => x"38811977",
   250 => x"812a5859",
   251 => x"76f738f7",
   252 => x"19769fff",
   253 => x"06545972",
   254 => x"802e8b38",
   255 => x"fc8016b6",
   256 => x"cc525698",
   257 => x"ad2d75b0",
   258 => x"80802e09",
   259 => x"81068938",
   260 => x"820bfedc",
   261 => x"0c88af04",
   262 => x"75988080",
   263 => x"2e098106",
   264 => x"8938810b",
   265 => x"fedc0c88",
   266 => x"af04800b",
   267 => x"fedc0c81",
   268 => x"5b807625",
   269 => x"80e93878",
   270 => x"52765184",
   271 => x"802db8b0",
   272 => x"52b6cc51",
   273 => x"98da2db6",
   274 => x"b008802e",
   275 => x"bb38b8b0",
   276 => x"5a83fc58",
   277 => x"79708405",
   278 => x"5b087083",
   279 => x"fe800671",
   280 => x"882b83fe",
   281 => x"80067188",
   282 => x"2a077288",
   283 => x"2a83fe80",
   284 => x"0673982a",
   285 => x"07fec80c",
   286 => x"fec80c56",
   287 => x"fc195953",
   288 => x"778025d0",
   289 => x"38898f04",
   290 => x"b6b0085b",
   291 => x"848056b6",
   292 => x"cc5198ad",
   293 => x"2dfc8016",
   294 => x"81185856",
   295 => x"88b1047a",
   296 => x"5372b6b0",
   297 => x"0c02ac05",
   298 => x"0d0402fc",
   299 => x"050da5ee",
   300 => x"2dfec451",
   301 => x"81710c82",
   302 => x"710c0284",
   303 => x"050d0402",
   304 => x"f4050d74",
   305 => x"10157084",
   306 => x"29b4b005",
   307 => x"70085551",
   308 => x"5272802e",
   309 => x"90387280",
   310 => x"f52d5271",
   311 => x"802e8638",
   312 => x"725187b4",
   313 => x"2db3a451",
   314 => x"a7cc2da5",
   315 => x"ee2d8051",
   316 => x"84e52d02",
   317 => x"8c050d04",
   318 => x"02e8050d",
   319 => x"80705656",
   320 => x"75b5e008",
   321 => x"25af38bc",
   322 => x"bc08762e",
   323 => x"a8387451",
   324 => x"95cf2db6",
   325 => x"b0080981",
   326 => x"0570b6b0",
   327 => x"08079f2a",
   328 => x"77058117",
   329 => x"57575275",
   330 => x"b5e00825",
   331 => x"8838bcbc",
   332 => x"087526da",
   333 => x"38805674",
   334 => x"bcbc0827",
   335 => x"80d03874",
   336 => x"5195cf2d",
   337 => x"75842b52",
   338 => x"b6b00880",
   339 => x"2eae38b6",
   340 => x"e0128117",
   341 => x"b6b00856",
   342 => x"57528a53",
   343 => x"73708105",
   344 => x"5580f52d",
   345 => x"72708105",
   346 => x"5481b72d",
   347 => x"ff135372",
   348 => x"8025e938",
   349 => x"807281b7",
   350 => x"2d8b8504",
   351 => x"b6b008b6",
   352 => x"e01381b7",
   353 => x"2d811555",
   354 => x"8b7625ff",
   355 => x"aa380298",
   356 => x"050d0402",
   357 => x"fc050d72",
   358 => x"5170fd2e",
   359 => x"ad3870fd",
   360 => x"248a3870",
   361 => x"fc2e80c4",
   362 => x"388bf404",
   363 => x"70fe2eb1",
   364 => x"3870ff2e",
   365 => x"098106bc",
   366 => x"38b5e008",
   367 => x"5170802e",
   368 => x"b338ff11",
   369 => x"b5e00c8b",
   370 => x"f404b5e0",
   371 => x"08f00570",
   372 => x"b5e00c51",
   373 => x"7080259c",
   374 => x"38800bb5",
   375 => x"e00c8bf4",
   376 => x"04b5e008",
   377 => x"8105b5e0",
   378 => x"0c8bf404",
   379 => x"b5e00890",
   380 => x"05b5e00c",
   381 => x"89f82da6",
   382 => x"b12d0284",
   383 => x"050d0402",
   384 => x"fc050db6",
   385 => x"d808fb06",
   386 => x"b6d80c72",
   387 => x"5189bf2d",
   388 => x"0284050d",
   389 => x"0402fc05",
   390 => x"0db6d808",
   391 => x"8407b6d8",
   392 => x"0c725189",
   393 => x"bf2d0284",
   394 => x"050d0402",
   395 => x"fc050d80",
   396 => x"0bb5e00c",
   397 => x"89f82db4",
   398 => x"ac51a7cc",
   399 => x"2db49451",
   400 => x"a7dc2d02",
   401 => x"84050d04",
   402 => x"02f8050d",
   403 => x"bd900882",
   404 => x"06b3c40b",
   405 => x"80f52d52",
   406 => x"5270802e",
   407 => x"85387181",
   408 => x"0752b3dc",
   409 => x"0b80f52d",
   410 => x"5170802e",
   411 => x"85387184",
   412 => x"0752b6dc",
   413 => x"08802e85",
   414 => x"38719007",
   415 => x"5271b6b0",
   416 => x"0c028805",
   417 => x"0d0402f4",
   418 => x"050d810b",
   419 => x"b6dc0c90",
   420 => x"5186922d",
   421 => x"810bfec4",
   422 => x"0c900bfe",
   423 => x"c00c840b",
   424 => x"fec40c83",
   425 => x"0bfecc0c",
   426 => x"a3bc2da5",
   427 => x"cf2da3a1",
   428 => x"2da3a12d",
   429 => x"81f72d81",
   430 => x"5184e52d",
   431 => x"a3a12da3",
   432 => x"a12d8151",
   433 => x"84e52db1",
   434 => x"c45185f1",
   435 => x"2d84529d",
   436 => x"b32d8fbd",
   437 => x"2db6b008",
   438 => x"802e8638",
   439 => x"fe528de9",
   440 => x"04ff1252",
   441 => x"718024e7",
   442 => x"3871802e",
   443 => x"81813886",
   444 => x"c22db1dc",
   445 => x"5187b42d",
   446 => x"b6b00880",
   447 => x"2e8f38b3",
   448 => x"a451a7cc",
   449 => x"2d805184",
   450 => x"e52d8e97",
   451 => x"04b6b008",
   452 => x"518cab2d",
   453 => x"a5db2da3",
   454 => x"d42da7e1",
   455 => x"2db6b008",
   456 => x"bd940888",
   457 => x"2bbd9808",
   458 => x"07fed80c",
   459 => x"538cc82d",
   460 => x"b6b008b6",
   461 => x"d8082ea2",
   462 => x"38b6b008",
   463 => x"b6d80cb6",
   464 => x"b008fec0",
   465 => x"0c845272",
   466 => x"5184e52d",
   467 => x"a3a12da3",
   468 => x"a12dff12",
   469 => x"52718025",
   470 => x"ee387280",
   471 => x"2e89388a",
   472 => x"0bfec40c",
   473 => x"8e970482",
   474 => x"0bfec40c",
   475 => x"8e9704b1",
   476 => x"e85185f1",
   477 => x"2d800bb6",
   478 => x"b00c028c",
   479 => x"050d0402",
   480 => x"e8050d77",
   481 => x"797b5855",
   482 => x"55805372",
   483 => x"7625a338",
   484 => x"74708105",
   485 => x"5680f52d",
   486 => x"74708105",
   487 => x"5680f52d",
   488 => x"52527171",
   489 => x"2e863881",
   490 => x"518fb404",
   491 => x"8113538f",
   492 => x"8b048051",
   493 => x"70b6b00c",
   494 => x"0298050d",
   495 => x"0402d805",
   496 => x"0d800bbc",
   497 => x"b80cb8b0",
   498 => x"528051a0",
   499 => x"9b2db6b0",
   500 => x"0854b6b0",
   501 => x"088c38b1",
   502 => x"fc5185f1",
   503 => x"2d735594",
   504 => x"d8048056",
   505 => x"810bbcdc",
   506 => x"0c8853b2",
   507 => x"8852b8e6",
   508 => x"518eff2d",
   509 => x"b6b00876",
   510 => x"2e098106",
   511 => x"8738b6b0",
   512 => x"08bcdc0c",
   513 => x"8853b294",
   514 => x"52b98251",
   515 => x"8eff2db6",
   516 => x"b0088738",
   517 => x"b6b008bc",
   518 => x"dc0cbcdc",
   519 => x"08802e80",
   520 => x"f638bbf6",
   521 => x"0b80f52d",
   522 => x"bbf70b80",
   523 => x"f52d7198",
   524 => x"2b71902b",
   525 => x"07bbf80b",
   526 => x"80f52d70",
   527 => x"882b7207",
   528 => x"bbf90b80",
   529 => x"f52d7107",
   530 => x"bcae0b80",
   531 => x"f52dbcaf",
   532 => x"0b80f52d",
   533 => x"71882b07",
   534 => x"535f5452",
   535 => x"5a565755",
   536 => x"7381abaa",
   537 => x"2e098106",
   538 => x"8d387551",
   539 => x"a1bb2db6",
   540 => x"b0085691",
   541 => x"83047382",
   542 => x"d4d52e87",
   543 => x"38b2a051",
   544 => x"91c404b8",
   545 => x"b0527551",
   546 => x"a09b2db6",
   547 => x"b00855b6",
   548 => x"b008802e",
   549 => x"83c23888",
   550 => x"53b29452",
   551 => x"b982518e",
   552 => x"ff2db6b0",
   553 => x"08893881",
   554 => x"0bbcb80c",
   555 => x"91ca0488",
   556 => x"53b28852",
   557 => x"b8e6518e",
   558 => x"ff2db6b0",
   559 => x"08802e8a",
   560 => x"38b2b451",
   561 => x"85f12d92",
   562 => x"a404bcae",
   563 => x"0b80f52d",
   564 => x"547380d5",
   565 => x"2e098106",
   566 => x"80ca38bc",
   567 => x"af0b80f5",
   568 => x"2d547381",
   569 => x"aa2e0981",
   570 => x"06ba3880",
   571 => x"0bb8b00b",
   572 => x"80f52d56",
   573 => x"547481e9",
   574 => x"2e833881",
   575 => x"547481eb",
   576 => x"2e8c3880",
   577 => x"5573752e",
   578 => x"09810682",
   579 => x"cb38b8bb",
   580 => x"0b80f52d",
   581 => x"55748d38",
   582 => x"b8bc0b80",
   583 => x"f52d5473",
   584 => x"822e8638",
   585 => x"805594d8",
   586 => x"04b8bd0b",
   587 => x"80f52d70",
   588 => x"bcb00cff",
   589 => x"05bcb40c",
   590 => x"b8be0b80",
   591 => x"f52db8bf",
   592 => x"0b80f52d",
   593 => x"58760577",
   594 => x"82802905",
   595 => x"70bcc00c",
   596 => x"b8c00b80",
   597 => x"f52d70bc",
   598 => x"d40cbcb8",
   599 => x"08595758",
   600 => x"76802e81",
   601 => x"a3388853",
   602 => x"b29452b9",
   603 => x"82518eff",
   604 => x"2db6b008",
   605 => x"81e238bc",
   606 => x"b0087084",
   607 => x"2bbcbc0c",
   608 => x"70bcd00c",
   609 => x"b8d50b80",
   610 => x"f52db8d4",
   611 => x"0b80f52d",
   612 => x"71828029",
   613 => x"05b8d60b",
   614 => x"80f52d70",
   615 => x"84808029",
   616 => x"12b8d70b",
   617 => x"80f52d70",
   618 => x"81800a29",
   619 => x"1270bcd8",
   620 => x"0cbcd408",
   621 => x"7129bcc0",
   622 => x"080570bc",
   623 => x"c40cb8dd",
   624 => x"0b80f52d",
   625 => x"b8dc0b80",
   626 => x"f52d7182",
   627 => x"802905b8",
   628 => x"de0b80f5",
   629 => x"2d708480",
   630 => x"802912b8",
   631 => x"df0b80f5",
   632 => x"2d70982b",
   633 => x"81f00a06",
   634 => x"720570bc",
   635 => x"c80cfe11",
   636 => x"7e297705",
   637 => x"bccc0c52",
   638 => x"59524354",
   639 => x"5e515259",
   640 => x"525d5759",
   641 => x"5794d604",
   642 => x"b8c20b80",
   643 => x"f52db8c1",
   644 => x"0b80f52d",
   645 => x"71828029",
   646 => x"0570bcbc",
   647 => x"0c70a029",
   648 => x"83ff0570",
   649 => x"892a70bc",
   650 => x"d00cb8c7",
   651 => x"0b80f52d",
   652 => x"b8c60b80",
   653 => x"f52d7182",
   654 => x"80290570",
   655 => x"bcd80c7b",
   656 => x"71291e70",
   657 => x"bccc0c7d",
   658 => x"bcc80c73",
   659 => x"05bcc40c",
   660 => x"555e5151",
   661 => x"55558155",
   662 => x"74b6b00c",
   663 => x"02a8050d",
   664 => x"0402ec05",
   665 => x"0d767087",
   666 => x"2c7180ff",
   667 => x"06555654",
   668 => x"bcb8088a",
   669 => x"3873882c",
   670 => x"7481ff06",
   671 => x"5455b8b0",
   672 => x"52bcc008",
   673 => x"1551a09b",
   674 => x"2db6b008",
   675 => x"54b6b008",
   676 => x"802eb338",
   677 => x"bcb80880",
   678 => x"2e983872",
   679 => x"8429b8b0",
   680 => x"05700852",
   681 => x"53a1bb2d",
   682 => x"b6b008f0",
   683 => x"0a065395",
   684 => x"c4047210",
   685 => x"b8b00570",
   686 => x"80e02d52",
   687 => x"53a1eb2d",
   688 => x"b6b00853",
   689 => x"725473b6",
   690 => x"b00c0294",
   691 => x"050d0402",
   692 => x"ec050d76",
   693 => x"70842cbc",
   694 => x"cc080571",
   695 => x"8f065255",
   696 => x"53728938",
   697 => x"b8b05273",
   698 => x"51a09b2d",
   699 => x"72a029b8",
   700 => x"b0055480",
   701 => x"7480f52d",
   702 => x"54557275",
   703 => x"2e833881",
   704 => x"557281e5",
   705 => x"2e933874",
   706 => x"802e8e38",
   707 => x"8b1480f5",
   708 => x"2d980653",
   709 => x"72802e83",
   710 => x"38805473",
   711 => x"b6b00c02",
   712 => x"94050d04",
   713 => x"02cc050d",
   714 => x"7e605e5a",
   715 => x"800bbcc8",
   716 => x"08bccc08",
   717 => x"595c5680",
   718 => x"58bcbc08",
   719 => x"782e81ae",
   720 => x"38778f06",
   721 => x"a0175754",
   722 => x"738f38b8",
   723 => x"b0527651",
   724 => x"811757a0",
   725 => x"9b2db8b0",
   726 => x"56807680",
   727 => x"f52d5654",
   728 => x"74742e83",
   729 => x"38815474",
   730 => x"81e52e80",
   731 => x"f6388170",
   732 => x"7506555c",
   733 => x"73802e80",
   734 => x"ea388b16",
   735 => x"80f52d98",
   736 => x"06597880",
   737 => x"de388b53",
   738 => x"7c527551",
   739 => x"8eff2db6",
   740 => x"b00880cf",
   741 => x"389c1608",
   742 => x"51a1bb2d",
   743 => x"b6b00884",
   744 => x"1b0c9a16",
   745 => x"80e02d51",
   746 => x"a1eb2db6",
   747 => x"b008b6b0",
   748 => x"08881c0c",
   749 => x"b6b00855",
   750 => x"55bcb808",
   751 => x"802e9838",
   752 => x"941680e0",
   753 => x"2d51a1eb",
   754 => x"2db6b008",
   755 => x"902b83ff",
   756 => x"f00a0670",
   757 => x"16515473",
   758 => x"881b0c78",
   759 => x"7a0c7b54",
   760 => x"98a40481",
   761 => x"1858bcbc",
   762 => x"087826fe",
   763 => x"d438bcb8",
   764 => x"08802eae",
   765 => x"387a5194",
   766 => x"e12db6b0",
   767 => x"08b6b008",
   768 => x"80ffffff",
   769 => x"f806555b",
   770 => x"7380ffff",
   771 => x"fff82e92",
   772 => x"38b6b008",
   773 => x"fe05bcb0",
   774 => x"0829bcc4",
   775 => x"08055796",
   776 => x"b7048054",
   777 => x"73b6b00c",
   778 => x"02b4050d",
   779 => x"0402f405",
   780 => x"0d747008",
   781 => x"8105710c",
   782 => x"7008bcb4",
   783 => x"08065353",
   784 => x"718e3888",
   785 => x"13085194",
   786 => x"e12db6b0",
   787 => x"0888140c",
   788 => x"810bb6b0",
   789 => x"0c028c05",
   790 => x"0d0402f0",
   791 => x"050d7588",
   792 => x"1108fe05",
   793 => x"bcb00829",
   794 => x"bcc40811",
   795 => x"7208bcb4",
   796 => x"08060579",
   797 => x"55535454",
   798 => x"a09b2d02",
   799 => x"90050d04",
   800 => x"02f0050d",
   801 => x"75881108",
   802 => x"fe05bcb0",
   803 => x"0829bcc4",
   804 => x"08117208",
   805 => x"bcb40806",
   806 => x"05795553",
   807 => x"54549edb",
   808 => x"2d029005",
   809 => x"0d0402f4",
   810 => x"050dd452",
   811 => x"81ff720c",
   812 => x"71085381",
   813 => x"ff720c72",
   814 => x"882b83fe",
   815 => x"80067208",
   816 => x"7081ff06",
   817 => x"51525381",
   818 => x"ff720c72",
   819 => x"7107882b",
   820 => x"72087081",
   821 => x"ff065152",
   822 => x"5381ff72",
   823 => x"0c727107",
   824 => x"882b7208",
   825 => x"7081ff06",
   826 => x"7207b6b0",
   827 => x"0c525302",
   828 => x"8c050d04",
   829 => x"02f4050d",
   830 => x"74767181",
   831 => x"ff06d40c",
   832 => x"5353bce0",
   833 => x"08853871",
   834 => x"892b5271",
   835 => x"982ad40c",
   836 => x"71902a70",
   837 => x"81ff06d4",
   838 => x"0c517188",
   839 => x"2a7081ff",
   840 => x"06d40c51",
   841 => x"7181ff06",
   842 => x"d40c7290",
   843 => x"2a7081ff",
   844 => x"06d40c51",
   845 => x"d4087081",
   846 => x"ff065151",
   847 => x"82b8bf52",
   848 => x"7081ff2e",
   849 => x"09810694",
   850 => x"3881ff0b",
   851 => x"d40cd408",
   852 => x"7081ff06",
   853 => x"ff145451",
   854 => x"5171e538",
   855 => x"70b6b00c",
   856 => x"028c050d",
   857 => x"0402fc05",
   858 => x"0d81c751",
   859 => x"81ff0bd4",
   860 => x"0cff1151",
   861 => x"708025f4",
   862 => x"38028405",
   863 => x"0d0402f0",
   864 => x"050d9ae5",
   865 => x"2d8fcf53",
   866 => x"805287fc",
   867 => x"80f75199",
   868 => x"f42db6b0",
   869 => x"0854b6b0",
   870 => x"08812e09",
   871 => x"8106a338",
   872 => x"81ff0bd4",
   873 => x"0c820a52",
   874 => x"849c80e9",
   875 => x"5199f42d",
   876 => x"b6b0088b",
   877 => x"3881ff0b",
   878 => x"d40c7353",
   879 => x"9bc8049a",
   880 => x"e52dff13",
   881 => x"5372c138",
   882 => x"72b6b00c",
   883 => x"0290050d",
   884 => x"0402f405",
   885 => x"0d81ff0b",
   886 => x"d40c9353",
   887 => x"805287fc",
   888 => x"80c15199",
   889 => x"f42db6b0",
   890 => x"088b3881",
   891 => x"ff0bd40c",
   892 => x"81539bfe",
   893 => x"049ae52d",
   894 => x"ff135372",
   895 => x"df3872b6",
   896 => x"b00c028c",
   897 => x"050d0402",
   898 => x"f0050d9a",
   899 => x"e52d83aa",
   900 => x"52849c80",
   901 => x"c85199f4",
   902 => x"2db6b008",
   903 => x"812e0981",
   904 => x"06923899",
   905 => x"a62db6b0",
   906 => x"0883ffff",
   907 => x"06537283",
   908 => x"aa2e9738",
   909 => x"9bd12d9c",
   910 => x"c5048154",
   911 => x"9daa04b2",
   912 => x"c05185f1",
   913 => x"2d80549d",
   914 => x"aa0481ff",
   915 => x"0bd40cb1",
   916 => x"539afe2d",
   917 => x"b6b00880",
   918 => x"2e80c038",
   919 => x"805287fc",
   920 => x"80fa5199",
   921 => x"f42db6b0",
   922 => x"08b13881",
   923 => x"ff0bd40c",
   924 => x"d4085381",
   925 => x"ff0bd40c",
   926 => x"81ff0bd4",
   927 => x"0c81ff0b",
   928 => x"d40c81ff",
   929 => x"0bd40c72",
   930 => x"862a7081",
   931 => x"06b6b008",
   932 => x"56515372",
   933 => x"802e9338",
   934 => x"9cba0472",
   935 => x"822eff9f",
   936 => x"38ff1353",
   937 => x"72ffaa38",
   938 => x"725473b6",
   939 => x"b00c0290",
   940 => x"050d0402",
   941 => x"f0050d81",
   942 => x"0bbce00c",
   943 => x"8454d008",
   944 => x"708f2a70",
   945 => x"81065151",
   946 => x"5372f338",
   947 => x"72d00c9a",
   948 => x"e52db2d0",
   949 => x"5185f12d",
   950 => x"d008708f",
   951 => x"2a708106",
   952 => x"51515372",
   953 => x"f338810b",
   954 => x"d00cb153",
   955 => x"805284d4",
   956 => x"80c05199",
   957 => x"f42db6b0",
   958 => x"08812ea1",
   959 => x"3872822e",
   960 => x"0981068c",
   961 => x"38b2dc51",
   962 => x"85f12d80",
   963 => x"539ed204",
   964 => x"ff135372",
   965 => x"d738ff14",
   966 => x"5473ffa2",
   967 => x"389c872d",
   968 => x"b6b008bc",
   969 => x"e00cb6b0",
   970 => x"088b3881",
   971 => x"5287fc80",
   972 => x"d05199f4",
   973 => x"2d81ff0b",
   974 => x"d40cd008",
   975 => x"708f2a70",
   976 => x"81065151",
   977 => x"5372f338",
   978 => x"72d00c81",
   979 => x"ff0bd40c",
   980 => x"815372b6",
   981 => x"b00c0290",
   982 => x"050d0402",
   983 => x"e8050d78",
   984 => x"5681ff0b",
   985 => x"d40cd008",
   986 => x"708f2a70",
   987 => x"81065151",
   988 => x"5372f338",
   989 => x"82810bd0",
   990 => x"0c81ff0b",
   991 => x"d40c7752",
   992 => x"87fc80d8",
   993 => x"5199f42d",
   994 => x"b6b00880",
   995 => x"2e8c38b2",
   996 => x"f45185f1",
   997 => x"2d8153a0",
   998 => x"920481ff",
   999 => x"0bd40c81",
  1000 => x"fe0bd40c",
  1001 => x"80ff5575",
  1002 => x"70840557",
  1003 => x"0870982a",
  1004 => x"d40c7090",
  1005 => x"2c7081ff",
  1006 => x"06d40c54",
  1007 => x"70882c70",
  1008 => x"81ff06d4",
  1009 => x"0c547081",
  1010 => x"ff06d40c",
  1011 => x"54ff1555",
  1012 => x"748025d3",
  1013 => x"3881ff0b",
  1014 => x"d40c81ff",
  1015 => x"0bd40c81",
  1016 => x"ff0bd40c",
  1017 => x"868da054",
  1018 => x"81ff0bd4",
  1019 => x"0cd40881",
  1020 => x"ff065574",
  1021 => x"8738ff14",
  1022 => x"5473ed38",
  1023 => x"81ff0bd4",
  1024 => x"0cd00870",
  1025 => x"8f2a7081",
  1026 => x"06515153",
  1027 => x"72f33872",
  1028 => x"d00c72b6",
  1029 => x"b00c0298",
  1030 => x"050d0402",
  1031 => x"e8050d78",
  1032 => x"55805681",
  1033 => x"ff0bd40c",
  1034 => x"d008708f",
  1035 => x"2a708106",
  1036 => x"51515372",
  1037 => x"f3388281",
  1038 => x"0bd00c81",
  1039 => x"ff0bd40c",
  1040 => x"775287fc",
  1041 => x"80d15199",
  1042 => x"f42d80db",
  1043 => x"c6df54b6",
  1044 => x"b008802e",
  1045 => x"8a38b384",
  1046 => x"5185f12d",
  1047 => x"a1b20481",
  1048 => x"ff0bd40c",
  1049 => x"d4087081",
  1050 => x"ff065153",
  1051 => x"7281fe2e",
  1052 => x"0981069d",
  1053 => x"3880ff53",
  1054 => x"99a62db6",
  1055 => x"b0087570",
  1056 => x"8405570c",
  1057 => x"ff135372",
  1058 => x"8025ed38",
  1059 => x"8156a197",
  1060 => x"04ff1454",
  1061 => x"73c93881",
  1062 => x"ff0bd40c",
  1063 => x"81ff0bd4",
  1064 => x"0cd00870",
  1065 => x"8f2a7081",
  1066 => x"06515153",
  1067 => x"72f33872",
  1068 => x"d00c75b6",
  1069 => x"b00c0298",
  1070 => x"050d0402",
  1071 => x"f4050d74",
  1072 => x"70882a83",
  1073 => x"fe800670",
  1074 => x"72982a07",
  1075 => x"72882b87",
  1076 => x"fc808006",
  1077 => x"73982b81",
  1078 => x"f00a0671",
  1079 => x"730707b6",
  1080 => x"b00c5651",
  1081 => x"5351028c",
  1082 => x"050d0402",
  1083 => x"f8050d02",
  1084 => x"8e0580f5",
  1085 => x"2d74882b",
  1086 => x"077083ff",
  1087 => x"ff06b6b0",
  1088 => x"0c510288",
  1089 => x"050d0402",
  1090 => x"fc050d72",
  1091 => x"5180710c",
  1092 => x"800b8412",
  1093 => x"0c028405",
  1094 => x"0d0402f0",
  1095 => x"050d7570",
  1096 => x"08841208",
  1097 => x"535353ff",
  1098 => x"5471712e",
  1099 => x"a838a5d5",
  1100 => x"2d841308",
  1101 => x"70842914",
  1102 => x"88117008",
  1103 => x"7081ff06",
  1104 => x"84180881",
  1105 => x"11870684",
  1106 => x"1a0c5351",
  1107 => x"55515151",
  1108 => x"a5cf2d71",
  1109 => x"5473b6b0",
  1110 => x"0c029005",
  1111 => x"0d0402f8",
  1112 => x"050da5d5",
  1113 => x"2de00870",
  1114 => x"8b2a7081",
  1115 => x"06515252",
  1116 => x"70802e9d",
  1117 => x"38bce408",
  1118 => x"708429bc",
  1119 => x"ec057381",
  1120 => x"ff06710c",
  1121 => x"5151bce4",
  1122 => x"08811187",
  1123 => x"06bce40c",
  1124 => x"51800bbd",
  1125 => x"8c0ca5c8",
  1126 => x"2da5cf2d",
  1127 => x"0288050d",
  1128 => x"0402fc05",
  1129 => x"0da5d52d",
  1130 => x"810bbd8c",
  1131 => x"0ca5cf2d",
  1132 => x"bd8c0851",
  1133 => x"70fa3802",
  1134 => x"84050d04",
  1135 => x"02fc050d",
  1136 => x"bce451a2",
  1137 => x"872da2de",
  1138 => x"51a5c42d",
  1139 => x"a4ee2d02",
  1140 => x"84050d04",
  1141 => x"02f4050d",
  1142 => x"a4d604b6",
  1143 => x"b00881f0",
  1144 => x"2e098106",
  1145 => x"8938810b",
  1146 => x"b6a40ca4",
  1147 => x"d604b6b0",
  1148 => x"0881e02e",
  1149 => x"09810689",
  1150 => x"38810bb6",
  1151 => x"a80ca4d6",
  1152 => x"04b6b008",
  1153 => x"52b6a808",
  1154 => x"802e8838",
  1155 => x"b6b00881",
  1156 => x"80055271",
  1157 => x"842c728f",
  1158 => x"065353b6",
  1159 => x"a408802e",
  1160 => x"99387284",
  1161 => x"29b5e405",
  1162 => x"72138171",
  1163 => x"2b700973",
  1164 => x"0806730c",
  1165 => x"515353a4",
  1166 => x"cc047284",
  1167 => x"29b5e405",
  1168 => x"72138371",
  1169 => x"2b720807",
  1170 => x"720c5353",
  1171 => x"800bb6a8",
  1172 => x"0c800bb6",
  1173 => x"a40cbce4",
  1174 => x"51a29a2d",
  1175 => x"b6b008ff",
  1176 => x"24fef838",
  1177 => x"800bb6b0",
  1178 => x"0c028c05",
  1179 => x"0d0402f8",
  1180 => x"050db5e4",
  1181 => x"528f5180",
  1182 => x"72708405",
  1183 => x"540cff11",
  1184 => x"51708025",
  1185 => x"f2380288",
  1186 => x"050d0402",
  1187 => x"f0050d75",
  1188 => x"51a5d52d",
  1189 => x"70822cfc",
  1190 => x"06b5e411",
  1191 => x"72109e06",
  1192 => x"71087072",
  1193 => x"2a708306",
  1194 => x"82742b70",
  1195 => x"09740676",
  1196 => x"0c545156",
  1197 => x"57535153",
  1198 => x"a5cf2d71",
  1199 => x"b6b00c02",
  1200 => x"90050d04",
  1201 => x"71980c04",
  1202 => x"ffb008b6",
  1203 => x"b00c0481",
  1204 => x"0bffb00c",
  1205 => x"04800bff",
  1206 => x"b00c0402",
  1207 => x"fc050d81",
  1208 => x"0bb6ac0c",
  1209 => x"815184e5",
  1210 => x"2d028405",
  1211 => x"0d0402fc",
  1212 => x"050d800b",
  1213 => x"b6ac0c80",
  1214 => x"5184e52d",
  1215 => x"0284050d",
  1216 => x"0402ec05",
  1217 => x"0d765480",
  1218 => x"52870b88",
  1219 => x"1580f52d",
  1220 => x"56537472",
  1221 => x"248338a0",
  1222 => x"53725182",
  1223 => x"ee2d8112",
  1224 => x"8b1580f5",
  1225 => x"2d545272",
  1226 => x"7225de38",
  1227 => x"0294050d",
  1228 => x"0402f005",
  1229 => x"0dbd9c08",
  1230 => x"5481f72d",
  1231 => x"800bbda0",
  1232 => x"0c730880",
  1233 => x"2e818038",
  1234 => x"820bb6c4",
  1235 => x"0cbda008",
  1236 => x"8f06b6c0",
  1237 => x"0c730852",
  1238 => x"71832e96",
  1239 => x"38718326",
  1240 => x"89387181",
  1241 => x"2eaf38a7",
  1242 => x"b2047185",
  1243 => x"2e9f38a7",
  1244 => x"b2048814",
  1245 => x"80f52d84",
  1246 => x"1508b394",
  1247 => x"53545285",
  1248 => x"f12d7184",
  1249 => x"29137008",
  1250 => x"5252a7b6",
  1251 => x"047351a6",
  1252 => x"812da7b2",
  1253 => x"04bd9008",
  1254 => x"8815082c",
  1255 => x"70810651",
  1256 => x"5271802e",
  1257 => x"8738b398",
  1258 => x"51a7af04",
  1259 => x"b39c5185",
  1260 => x"f12d8414",
  1261 => x"085185f1",
  1262 => x"2dbda008",
  1263 => x"8105bda0",
  1264 => x"0c8c1454",
  1265 => x"a6c10402",
  1266 => x"90050d04",
  1267 => x"71bd9c0c",
  1268 => x"a6b12dbd",
  1269 => x"a008ff05",
  1270 => x"bda40c04",
  1271 => x"71bda80c",
  1272 => x"0402e805",
  1273 => x"0dbd9c08",
  1274 => x"bda80857",
  1275 => x"5580f851",
  1276 => x"a58b2db6",
  1277 => x"b008812a",
  1278 => x"70810651",
  1279 => x"52719b38",
  1280 => x"8751a58b",
  1281 => x"2db6b008",
  1282 => x"812a7081",
  1283 => x"06515271",
  1284 => x"802eb138",
  1285 => x"a89a04a3",
  1286 => x"d42d8751",
  1287 => x"a58b2db6",
  1288 => x"b008f438",
  1289 => x"a8aa04a3",
  1290 => x"d42d80f8",
  1291 => x"51a58b2d",
  1292 => x"b6b008f3",
  1293 => x"38b6ac08",
  1294 => x"813270b6",
  1295 => x"ac0c7052",
  1296 => x"5284e52d",
  1297 => x"800bbd94",
  1298 => x"0c800bbd",
  1299 => x"980cb6ac",
  1300 => x"0882dd38",
  1301 => x"80da51a5",
  1302 => x"8b2db6b0",
  1303 => x"08802e8a",
  1304 => x"38bd9408",
  1305 => x"818007bd",
  1306 => x"940c80d9",
  1307 => x"51a58b2d",
  1308 => x"b6b00880",
  1309 => x"2e8a38bd",
  1310 => x"940880c0",
  1311 => x"07bd940c",
  1312 => x"819451a5",
  1313 => x"8b2db6b0",
  1314 => x"08802e89",
  1315 => x"38bd9408",
  1316 => x"9007bd94",
  1317 => x"0c819151",
  1318 => x"a58b2db6",
  1319 => x"b008802e",
  1320 => x"8938bd94",
  1321 => x"08a007bd",
  1322 => x"940c81f5",
  1323 => x"51a58b2d",
  1324 => x"b6b00880",
  1325 => x"2e8938bd",
  1326 => x"94088107",
  1327 => x"bd940c81",
  1328 => x"f251a58b",
  1329 => x"2db6b008",
  1330 => x"802e8938",
  1331 => x"bd940882",
  1332 => x"07bd940c",
  1333 => x"81eb51a5",
  1334 => x"8b2db6b0",
  1335 => x"08802e89",
  1336 => x"38bd9408",
  1337 => x"8407bd94",
  1338 => x"0c81f451",
  1339 => x"a58b2db6",
  1340 => x"b008802e",
  1341 => x"8938bd94",
  1342 => x"088807bd",
  1343 => x"940c80d8",
  1344 => x"51a58b2d",
  1345 => x"b6b00880",
  1346 => x"2e8a38bd",
  1347 => x"98088180",
  1348 => x"07bd980c",
  1349 => x"9251a58b",
  1350 => x"2db6b008",
  1351 => x"802e8a38",
  1352 => x"bd980880",
  1353 => x"c007bd98",
  1354 => x"0c9451a5",
  1355 => x"8b2db6b0",
  1356 => x"08802e89",
  1357 => x"38bd9808",
  1358 => x"9007bd98",
  1359 => x"0c9151a5",
  1360 => x"8b2db6b0",
  1361 => x"08802e89",
  1362 => x"38bd9808",
  1363 => x"a007bd98",
  1364 => x"0c9d51a5",
  1365 => x"8b2db6b0",
  1366 => x"08802e89",
  1367 => x"38bd9808",
  1368 => x"8107bd98",
  1369 => x"0c9b51a5",
  1370 => x"8b2db6b0",
  1371 => x"08802e89",
  1372 => x"38bd9808",
  1373 => x"8207bd98",
  1374 => x"0c9c51a5",
  1375 => x"8b2db6b0",
  1376 => x"08802e89",
  1377 => x"38bd9808",
  1378 => x"8407bd98",
  1379 => x"0ca351a5",
  1380 => x"8b2db6b0",
  1381 => x"08802e89",
  1382 => x"38bd9808",
  1383 => x"8807bd98",
  1384 => x"0c81fd51",
  1385 => x"a58b2d81",
  1386 => x"fa51a58b",
  1387 => x"2db09504",
  1388 => x"81f551a5",
  1389 => x"8b2db6b0",
  1390 => x"08812a70",
  1391 => x"81065152",
  1392 => x"71802eaf",
  1393 => x"38bda408",
  1394 => x"5271802e",
  1395 => x"8938ff12",
  1396 => x"bda40cab",
  1397 => x"f304bda0",
  1398 => x"0810bda0",
  1399 => x"08057084",
  1400 => x"29165152",
  1401 => x"88120880",
  1402 => x"2e8938ff",
  1403 => x"51881208",
  1404 => x"52712d81",
  1405 => x"f251a58b",
  1406 => x"2db6b008",
  1407 => x"812a7081",
  1408 => x"06515271",
  1409 => x"802eb138",
  1410 => x"bda008ff",
  1411 => x"11bda408",
  1412 => x"56535373",
  1413 => x"72258938",
  1414 => x"8114bda4",
  1415 => x"0cacb804",
  1416 => x"72101370",
  1417 => x"84291651",
  1418 => x"52881208",
  1419 => x"802e8938",
  1420 => x"fe518812",
  1421 => x"0852712d",
  1422 => x"81fd51a5",
  1423 => x"8b2db6b0",
  1424 => x"08812a70",
  1425 => x"81065152",
  1426 => x"71802e86",
  1427 => x"38800bbd",
  1428 => x"a40c81fa",
  1429 => x"51a58b2d",
  1430 => x"b6b00881",
  1431 => x"2a708106",
  1432 => x"51527180",
  1433 => x"2e8938bd",
  1434 => x"a008ff05",
  1435 => x"bda40cbd",
  1436 => x"a4087053",
  1437 => x"5473802e",
  1438 => x"8a388c15",
  1439 => x"ff155555",
  1440 => x"acf50482",
  1441 => x"0bb6c40c",
  1442 => x"718f06b6",
  1443 => x"c00c81eb",
  1444 => x"51a58b2d",
  1445 => x"b6b00881",
  1446 => x"2a708106",
  1447 => x"51527180",
  1448 => x"2ead3874",
  1449 => x"08852e09",
  1450 => x"8106a438",
  1451 => x"881580f5",
  1452 => x"2dff0552",
  1453 => x"71881681",
  1454 => x"b72d7198",
  1455 => x"2b527180",
  1456 => x"25883880",
  1457 => x"0b881681",
  1458 => x"b72d7451",
  1459 => x"a6812d81",
  1460 => x"f451a58b",
  1461 => x"2db6b008",
  1462 => x"812a7081",
  1463 => x"06515271",
  1464 => x"802eb338",
  1465 => x"7408852e",
  1466 => x"098106aa",
  1467 => x"38881580",
  1468 => x"f52d8105",
  1469 => x"52718816",
  1470 => x"81b72d71",
  1471 => x"81ff068b",
  1472 => x"1680f52d",
  1473 => x"54527272",
  1474 => x"27873872",
  1475 => x"881681b7",
  1476 => x"2d7451a6",
  1477 => x"812d80da",
  1478 => x"51a58b2d",
  1479 => x"b6b00881",
  1480 => x"2a708106",
  1481 => x"51527180",
  1482 => x"2e81a638",
  1483 => x"bd9c08bd",
  1484 => x"a4085553",
  1485 => x"73802e8a",
  1486 => x"388c13ff",
  1487 => x"155553ae",
  1488 => x"b4047208",
  1489 => x"5271822e",
  1490 => x"a6387182",
  1491 => x"26893871",
  1492 => x"812ea938",
  1493 => x"afd10471",
  1494 => x"832eb138",
  1495 => x"71842e09",
  1496 => x"810680ed",
  1497 => x"38881308",
  1498 => x"51a7cc2d",
  1499 => x"afd104bd",
  1500 => x"a4085188",
  1501 => x"13085271",
  1502 => x"2dafd104",
  1503 => x"810b8814",
  1504 => x"082bbd90",
  1505 => x"0832bd90",
  1506 => x"0cafa704",
  1507 => x"881380f5",
  1508 => x"2d81058b",
  1509 => x"1480f52d",
  1510 => x"53547174",
  1511 => x"24833880",
  1512 => x"54738814",
  1513 => x"81b72da6",
  1514 => x"b12dafd1",
  1515 => x"04750880",
  1516 => x"2ea23875",
  1517 => x"0851a58b",
  1518 => x"2db6b008",
  1519 => x"81065271",
  1520 => x"802e8b38",
  1521 => x"bda40851",
  1522 => x"84160852",
  1523 => x"712d8816",
  1524 => x"5675da38",
  1525 => x"8054800b",
  1526 => x"b6c40c73",
  1527 => x"8f06b6c0",
  1528 => x"0ca05273",
  1529 => x"bda4082e",
  1530 => x"09810698",
  1531 => x"38bda008",
  1532 => x"ff057432",
  1533 => x"70098105",
  1534 => x"7072079f",
  1535 => x"2a917131",
  1536 => x"51515353",
  1537 => x"715182ee",
  1538 => x"2d811454",
  1539 => x"8e7425c6",
  1540 => x"38b6ac08",
  1541 => x"5271b6b0",
  1542 => x"0c029805",
  1543 => x"0d040000",
  1544 => x"00ffffff",
  1545 => x"ff00ffff",
  1546 => x"ffff00ff",
  1547 => x"ffffff00",
  1548 => x"52657365",
  1549 => x"74000000",
  1550 => x"53617665",
  1551 => x"20736574",
  1552 => x"74696e67",
  1553 => x"73000000",
  1554 => x"5363616e",
  1555 => x"6c696e65",
  1556 => x"73000000",
  1557 => x"4c6f6164",
  1558 => x"20524f4d",
  1559 => x"20100000",
  1560 => x"45786974",
  1561 => x"00000000",
  1562 => x"50432045",
  1563 => x"6e67696e",
  1564 => x"65206d6f",
  1565 => x"64650000",
  1566 => x"54757262",
  1567 => x"6f677261",
  1568 => x"66782031",
  1569 => x"36206d6f",
  1570 => x"64650000",
  1571 => x"56474120",
  1572 => x"2d203331",
  1573 => x"4b487a2c",
  1574 => x"20363048",
  1575 => x"7a000000",
  1576 => x"5456202d",
  1577 => x"20343830",
  1578 => x"692c2036",
  1579 => x"30487a00",
  1580 => x"4261636b",
  1581 => x"00000000",
  1582 => x"46504741",
  1583 => x"50434520",
  1584 => x"43464700",
  1585 => x"496e6974",
  1586 => x"69616c69",
  1587 => x"7a696e67",
  1588 => x"20534420",
  1589 => x"63617264",
  1590 => x"0a000000",
  1591 => x"424f4f54",
  1592 => x"20202020",
  1593 => x"50434500",
  1594 => x"43617264",
  1595 => x"20696e69",
  1596 => x"74206661",
  1597 => x"696c6564",
  1598 => x"0a000000",
  1599 => x"4d425220",
  1600 => x"6661696c",
  1601 => x"0a000000",
  1602 => x"46415431",
  1603 => x"36202020",
  1604 => x"00000000",
  1605 => x"46415433",
  1606 => x"32202020",
  1607 => x"00000000",
  1608 => x"4e6f2070",
  1609 => x"61727469",
  1610 => x"74696f6e",
  1611 => x"20736967",
  1612 => x"0a000000",
  1613 => x"42616420",
  1614 => x"70617274",
  1615 => x"0a000000",
  1616 => x"53444843",
  1617 => x"20657272",
  1618 => x"6f72210a",
  1619 => x"00000000",
  1620 => x"53442069",
  1621 => x"6e69742e",
  1622 => x"2e2e0a00",
  1623 => x"53442063",
  1624 => x"61726420",
  1625 => x"72657365",
  1626 => x"74206661",
  1627 => x"696c6564",
  1628 => x"210a0000",
  1629 => x"57726974",
  1630 => x"65206661",
  1631 => x"696c6564",
  1632 => x"0a000000",
  1633 => x"52656164",
  1634 => x"20666169",
  1635 => x"6c65640a",
  1636 => x"00000000",
  1637 => x"16200000",
  1638 => x"14200000",
  1639 => x"15200000",
  1640 => x"00000002",
  1641 => x"00000002",
  1642 => x"00001830",
  1643 => x"000004aa",
  1644 => x"00000002",
  1645 => x"00001838",
  1646 => x"00000377",
  1647 => x"00000003",
  1648 => x"00001a0c",
  1649 => x"00000002",
  1650 => x"00000001",
  1651 => x"00001848",
  1652 => x"00000001",
  1653 => x"00000003",
  1654 => x"00001a04",
  1655 => x"00000002",
  1656 => x"00000002",
  1657 => x"00001854",
  1658 => x"0000062b",
  1659 => x"00000002",
  1660 => x"00001860",
  1661 => x"000012ee",
  1662 => x"00000000",
  1663 => x"00000000",
  1664 => x"00000000",
  1665 => x"00001868",
  1666 => x"00001878",
  1667 => x"0000188c",
  1668 => x"000018a0",
  1669 => x"0000004d",
  1670 => x"000005ff",
  1671 => x"0000002c",
  1672 => x"00000615",
  1673 => x"00000000",
  1674 => x"00000000",
  1675 => x"00000002",
  1676 => x"00001b60",
  1677 => x"000004bf",
  1678 => x"00000002",
  1679 => x"00001b70",
  1680 => x"000004bf",
  1681 => x"00000002",
  1682 => x"00001b80",
  1683 => x"000004bf",
  1684 => x"00000002",
  1685 => x"00001b90",
  1686 => x"000004bf",
  1687 => x"00000002",
  1688 => x"00001ba0",
  1689 => x"000004bf",
  1690 => x"00000002",
  1691 => x"00001bb0",
  1692 => x"000004bf",
  1693 => x"00000002",
  1694 => x"00001bc0",
  1695 => x"000004bf",
  1696 => x"00000002",
  1697 => x"00001bd0",
  1698 => x"000004bf",
  1699 => x"00000002",
  1700 => x"00001be0",
  1701 => x"000004bf",
  1702 => x"00000002",
  1703 => x"00001bf0",
  1704 => x"000004bf",
  1705 => x"00000002",
  1706 => x"00001c00",
  1707 => x"000004bf",
  1708 => x"00000002",
  1709 => x"00001c10",
  1710 => x"000004bf",
  1711 => x"00000002",
  1712 => x"00001c20",
  1713 => x"000004bf",
  1714 => x"00000004",
  1715 => x"000018b0",
  1716 => x"000019a4",
  1717 => x"00000000",
  1718 => x"00000000",
  1719 => x"00000593",
  1720 => x"00000000",
  1721 => x"00000000",
  1722 => x"00000000",
  1723 => x"00000000",
  1724 => x"00000000",
  1725 => x"00000000",
  1726 => x"00000000",
  1727 => x"00000000",
  1728 => x"00000000",
  1729 => x"00000000",
  1730 => x"00000000",
  1731 => x"00000000",
  1732 => x"00000000",
  1733 => x"00000000",
  1734 => x"00000000",
  1735 => x"00000000",
  1736 => x"00000000",
  1737 => x"00000000",
  1738 => x"00000000",
  1739 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

